magic
tech gf180mcuD
magscale 1 5
timestamp 1702171133
<< nwell >>
rect 629 173440 279371 173872
rect 629 172656 279371 173088
rect 629 171872 279371 172304
rect 629 171088 279371 171520
rect 629 170304 279371 170736
rect 629 169520 279371 169952
rect 629 168736 279371 169168
rect 629 167952 279371 168384
rect 629 167168 279371 167600
rect 629 166384 279371 166816
rect 629 165600 279371 166032
rect 629 164816 279371 165248
rect 629 164032 279371 164464
rect 629 163248 279371 163680
rect 629 162464 279371 162896
rect 629 161680 279371 162112
rect 629 160896 279371 161328
rect 629 160112 279371 160544
rect 629 159328 279371 159760
rect 629 158544 279371 158976
rect 629 157760 279371 158192
rect 629 156976 279371 157408
rect 629 156192 279371 156624
rect 629 155408 279371 155840
rect 629 154624 279371 155056
rect 629 153840 279371 154272
rect 629 153056 279371 153488
rect 629 152272 279371 152704
rect 629 151488 279371 151920
rect 629 150704 279371 151136
rect 629 149920 279371 150352
rect 629 149136 279371 149568
rect 629 148352 279371 148784
rect 629 147568 279371 148000
rect 629 146784 279371 147216
rect 629 146000 279371 146432
rect 629 145216 279371 145648
rect 629 144432 279371 144864
rect 629 143648 279371 144080
rect 629 142864 279371 143296
rect 629 142080 279371 142512
rect 629 141296 279371 141728
rect 629 140512 279371 140944
rect 629 139728 279371 140160
rect 629 138944 279371 139376
rect 629 138160 279371 138592
rect 629 137376 279371 137808
rect 629 136592 279371 137024
rect 629 135808 279371 136240
rect 629 135024 279371 135456
rect 629 134240 279371 134672
rect 629 133456 279371 133888
rect 629 132672 279371 133104
rect 629 131888 279371 132320
rect 629 131104 279371 131536
rect 629 130320 279371 130752
rect 629 129536 279371 129968
rect 629 128752 279371 129184
rect 629 127968 279371 128400
rect 629 127184 279371 127616
rect 629 126400 279371 126832
rect 629 125616 279371 126048
rect 629 124832 279371 125264
rect 629 124048 279371 124480
rect 629 123264 279371 123696
rect 629 122480 279371 122912
rect 629 121696 279371 122128
rect 629 120912 279371 121344
rect 629 120128 279371 120560
rect 629 119344 279371 119776
rect 629 118560 279371 118992
rect 629 117776 279371 118208
rect 629 116992 279371 117424
rect 629 116208 279371 116640
rect 629 115424 279371 115856
rect 629 114640 279371 115072
rect 629 113856 279371 114288
rect 629 113072 279371 113504
rect 629 112288 279371 112720
rect 629 111504 279371 111936
rect 629 110720 279371 111152
rect 629 109936 279371 110368
rect 629 109152 279371 109584
rect 629 108368 279371 108800
rect 629 107584 279371 108016
rect 629 106800 279371 107232
rect 629 106016 279371 106448
rect 629 105232 279371 105664
rect 629 104448 279371 104880
rect 629 103664 279371 104096
rect 629 102880 279371 103312
rect 629 102096 279371 102528
rect 629 101312 279371 101744
rect 629 100528 279371 100960
rect 629 99744 279371 100176
rect 629 98960 279371 99392
rect 629 98176 279371 98608
rect 629 97392 279371 97824
rect 629 96608 279371 97040
rect 629 95824 279371 96256
rect 629 95040 279371 95472
rect 629 94256 279371 94688
rect 629 93472 279371 93904
rect 629 92688 279371 93120
rect 629 91904 279371 92336
rect 629 91120 279371 91552
rect 629 90336 279371 90768
rect 629 89552 279371 89984
rect 629 88768 279371 89200
rect 629 87984 279371 88416
rect 629 87200 279371 87632
rect 629 86416 279371 86848
rect 629 85632 279371 86064
rect 629 84848 279371 85280
rect 629 84064 279371 84496
rect 629 83280 279371 83712
rect 629 82496 279371 82928
rect 629 81712 279371 82144
rect 629 80928 279371 81360
rect 629 80144 279371 80576
rect 629 79360 279371 79792
rect 629 78576 279371 79008
rect 629 77792 279371 78224
rect 629 77008 279371 77440
rect 629 76224 279371 76656
rect 629 75440 279371 75872
rect 629 74656 279371 75088
rect 629 73872 279371 74304
rect 629 73088 279371 73520
rect 629 72304 279371 72736
rect 629 71520 279371 71952
rect 629 70736 279371 71168
rect 629 69952 279371 70384
rect 629 69168 279371 69600
rect 629 68384 279371 68816
rect 629 67600 279371 68032
rect 629 66816 279371 67248
rect 629 66032 279371 66464
rect 629 65248 279371 65680
rect 629 64464 279371 64896
rect 629 63680 279371 64112
rect 629 62896 279371 63328
rect 629 62112 279371 62544
rect 629 61328 279371 61760
rect 629 60544 279371 60976
rect 629 59760 279371 60192
rect 629 58976 279371 59408
rect 629 58192 279371 58624
rect 629 57408 279371 57840
rect 629 56624 279371 57056
rect 629 55840 279371 56272
rect 629 55056 279371 55488
rect 629 54272 279371 54704
rect 629 53488 279371 53920
rect 629 52704 279371 53136
rect 629 51920 279371 52352
rect 629 51136 279371 51568
rect 629 50352 279371 50784
rect 629 49568 279371 50000
rect 629 48784 279371 49216
rect 629 48000 279371 48432
rect 629 47216 279371 47648
rect 629 46432 279371 46864
rect 629 45648 279371 46080
rect 629 44864 279371 45296
rect 629 44080 279371 44512
rect 629 43296 279371 43728
rect 629 42512 279371 42944
rect 629 41728 279371 42160
rect 629 40944 279371 41376
rect 629 40160 279371 40592
rect 629 39376 279371 39808
rect 629 38592 279371 39024
rect 629 37808 279371 38240
rect 629 37024 279371 37456
rect 629 36240 279371 36672
rect 629 35456 279371 35888
rect 629 34672 279371 35104
rect 629 33888 279371 34320
rect 629 33104 279371 33536
rect 629 32320 279371 32752
rect 629 31536 279371 31968
rect 629 30752 279371 31184
rect 629 29968 279371 30400
rect 629 29184 279371 29616
rect 629 28400 279371 28832
rect 629 27616 279371 28048
rect 629 26832 279371 27264
rect 629 26048 279371 26480
rect 629 25264 279371 25696
rect 629 24480 279371 24912
rect 629 23696 279371 24128
rect 629 22912 279371 23344
rect 629 22128 279371 22560
rect 629 21344 279371 21776
rect 629 20560 279371 20992
rect 629 19776 279371 20208
rect 629 18992 279371 19424
rect 629 18208 279371 18640
rect 629 17424 279371 17856
rect 629 16640 279371 17072
rect 629 15856 279371 16288
rect 629 15072 279371 15504
rect 629 14288 279371 14720
rect 629 13504 279371 13936
rect 629 12720 279371 13152
rect 629 11936 279371 12368
rect 629 11152 279371 11584
rect 629 10368 279371 10800
rect 629 9584 279371 10016
rect 629 8800 279371 9232
rect 629 8016 279371 8448
rect 629 7232 279371 7664
rect 629 6448 279371 6880
rect 629 5664 279371 6096
rect 629 4880 279371 5312
rect 629 4096 279371 4528
rect 629 3312 279371 3744
rect 629 2528 279371 2960
rect 629 1744 279371 2176
<< pwell >>
rect 629 173872 279371 174091
rect 629 173088 279371 173440
rect 629 172304 279371 172656
rect 629 171520 279371 171872
rect 629 170736 279371 171088
rect 629 169952 279371 170304
rect 629 169168 279371 169520
rect 629 168384 279371 168736
rect 629 167600 279371 167952
rect 629 166816 279371 167168
rect 629 166032 279371 166384
rect 629 165248 279371 165600
rect 629 164464 279371 164816
rect 629 163680 279371 164032
rect 629 162896 279371 163248
rect 629 162112 279371 162464
rect 629 161328 279371 161680
rect 629 160544 279371 160896
rect 629 159760 279371 160112
rect 629 158976 279371 159328
rect 629 158192 279371 158544
rect 629 157408 279371 157760
rect 629 156624 279371 156976
rect 629 155840 279371 156192
rect 629 155056 279371 155408
rect 629 154272 279371 154624
rect 629 153488 279371 153840
rect 629 152704 279371 153056
rect 629 151920 279371 152272
rect 629 151136 279371 151488
rect 629 150352 279371 150704
rect 629 149568 279371 149920
rect 629 148784 279371 149136
rect 629 148000 279371 148352
rect 629 147216 279371 147568
rect 629 146432 279371 146784
rect 629 145648 279371 146000
rect 629 144864 279371 145216
rect 629 144080 279371 144432
rect 629 143296 279371 143648
rect 629 142512 279371 142864
rect 629 141728 279371 142080
rect 629 140944 279371 141296
rect 629 140160 279371 140512
rect 629 139376 279371 139728
rect 629 138592 279371 138944
rect 629 137808 279371 138160
rect 629 137024 279371 137376
rect 629 136240 279371 136592
rect 629 135456 279371 135808
rect 629 134672 279371 135024
rect 629 133888 279371 134240
rect 629 133104 279371 133456
rect 629 132320 279371 132672
rect 629 131536 279371 131888
rect 629 130752 279371 131104
rect 629 129968 279371 130320
rect 629 129184 279371 129536
rect 629 128400 279371 128752
rect 629 127616 279371 127968
rect 629 126832 279371 127184
rect 629 126048 279371 126400
rect 629 125264 279371 125616
rect 629 124480 279371 124832
rect 629 123696 279371 124048
rect 629 122912 279371 123264
rect 629 122128 279371 122480
rect 629 121344 279371 121696
rect 629 120560 279371 120912
rect 629 119776 279371 120128
rect 629 118992 279371 119344
rect 629 118208 279371 118560
rect 629 117424 279371 117776
rect 629 116640 279371 116992
rect 629 115856 279371 116208
rect 629 115072 279371 115424
rect 629 114288 279371 114640
rect 629 113504 279371 113856
rect 629 112720 279371 113072
rect 629 111936 279371 112288
rect 629 111152 279371 111504
rect 629 110368 279371 110720
rect 629 109584 279371 109936
rect 629 108800 279371 109152
rect 629 108016 279371 108368
rect 629 107232 279371 107584
rect 629 106448 279371 106800
rect 629 105664 279371 106016
rect 629 104880 279371 105232
rect 629 104096 279371 104448
rect 629 103312 279371 103664
rect 629 102528 279371 102880
rect 629 101744 279371 102096
rect 629 100960 279371 101312
rect 629 100176 279371 100528
rect 629 99392 279371 99744
rect 629 98608 279371 98960
rect 629 97824 279371 98176
rect 629 97040 279371 97392
rect 629 96256 279371 96608
rect 629 95472 279371 95824
rect 629 94688 279371 95040
rect 629 93904 279371 94256
rect 629 93120 279371 93472
rect 629 92336 279371 92688
rect 629 91552 279371 91904
rect 629 90768 279371 91120
rect 629 89984 279371 90336
rect 629 89200 279371 89552
rect 629 88416 279371 88768
rect 629 87632 279371 87984
rect 629 86848 279371 87200
rect 629 86064 279371 86416
rect 629 85280 279371 85632
rect 629 84496 279371 84848
rect 629 83712 279371 84064
rect 629 82928 279371 83280
rect 629 82144 279371 82496
rect 629 81360 279371 81712
rect 629 80576 279371 80928
rect 629 79792 279371 80144
rect 629 79008 279371 79360
rect 629 78224 279371 78576
rect 629 77440 279371 77792
rect 629 76656 279371 77008
rect 629 75872 279371 76224
rect 629 75088 279371 75440
rect 629 74304 279371 74656
rect 629 73520 279371 73872
rect 629 72736 279371 73088
rect 629 71952 279371 72304
rect 629 71168 279371 71520
rect 629 70384 279371 70736
rect 629 69600 279371 69952
rect 629 68816 279371 69168
rect 629 68032 279371 68384
rect 629 67248 279371 67600
rect 629 66464 279371 66816
rect 629 65680 279371 66032
rect 629 64896 279371 65248
rect 629 64112 279371 64464
rect 629 63328 279371 63680
rect 629 62544 279371 62896
rect 629 61760 279371 62112
rect 629 60976 279371 61328
rect 629 60192 279371 60544
rect 629 59408 279371 59760
rect 629 58624 279371 58976
rect 629 57840 279371 58192
rect 629 57056 279371 57408
rect 629 56272 279371 56624
rect 629 55488 279371 55840
rect 629 54704 279371 55056
rect 629 53920 279371 54272
rect 629 53136 279371 53488
rect 629 52352 279371 52704
rect 629 51568 279371 51920
rect 629 50784 279371 51136
rect 629 50000 279371 50352
rect 629 49216 279371 49568
rect 629 48432 279371 48784
rect 629 47648 279371 48000
rect 629 46864 279371 47216
rect 629 46080 279371 46432
rect 629 45296 279371 45648
rect 629 44512 279371 44864
rect 629 43728 279371 44080
rect 629 42944 279371 43296
rect 629 42160 279371 42512
rect 629 41376 279371 41728
rect 629 40592 279371 40944
rect 629 39808 279371 40160
rect 629 39024 279371 39376
rect 629 38240 279371 38592
rect 629 37456 279371 37808
rect 629 36672 279371 37024
rect 629 35888 279371 36240
rect 629 35104 279371 35456
rect 629 34320 279371 34672
rect 629 33536 279371 33888
rect 629 32752 279371 33104
rect 629 31968 279371 32320
rect 629 31184 279371 31536
rect 629 30400 279371 30752
rect 629 29616 279371 29968
rect 629 28832 279371 29184
rect 629 28048 279371 28400
rect 629 27264 279371 27616
rect 629 26480 279371 26832
rect 629 25696 279371 26048
rect 629 24912 279371 25264
rect 629 24128 279371 24480
rect 629 23344 279371 23696
rect 629 22560 279371 22912
rect 629 21776 279371 22128
rect 629 20992 279371 21344
rect 629 20208 279371 20560
rect 629 19424 279371 19776
rect 629 18640 279371 18992
rect 629 17856 279371 18208
rect 629 17072 279371 17424
rect 629 16288 279371 16640
rect 629 15504 279371 15856
rect 629 14720 279371 15072
rect 629 13936 279371 14288
rect 629 13152 279371 13504
rect 629 12368 279371 12720
rect 629 11584 279371 11936
rect 629 10800 279371 11152
rect 629 10016 279371 10368
rect 629 9232 279371 9584
rect 629 8448 279371 8800
rect 629 7664 279371 8016
rect 629 6880 279371 7232
rect 629 6096 279371 6448
rect 629 5312 279371 5664
rect 629 4528 279371 4880
rect 629 3744 279371 4096
rect 629 2960 279371 3312
rect 629 2176 279371 2528
rect 629 1525 279371 1744
<< obsm1 >>
rect 672 855 279328 174078
<< metal2 >>
rect 10192 0 10248 400
rect 11536 0 11592 400
rect 12880 0 12936 400
rect 14224 0 14280 400
rect 15568 0 15624 400
rect 16912 0 16968 400
rect 18256 0 18312 400
rect 19600 0 19656 400
rect 20944 0 21000 400
rect 22288 0 22344 400
rect 23632 0 23688 400
rect 24976 0 25032 400
rect 26320 0 26376 400
rect 27664 0 27720 400
rect 29008 0 29064 400
rect 30352 0 30408 400
rect 31696 0 31752 400
rect 33040 0 33096 400
rect 34384 0 34440 400
rect 35728 0 35784 400
rect 37072 0 37128 400
rect 38416 0 38472 400
rect 39760 0 39816 400
rect 41104 0 41160 400
rect 42448 0 42504 400
rect 43792 0 43848 400
rect 45136 0 45192 400
rect 46480 0 46536 400
rect 47824 0 47880 400
rect 49168 0 49224 400
rect 50512 0 50568 400
rect 51856 0 51912 400
rect 53200 0 53256 400
rect 54544 0 54600 400
rect 55888 0 55944 400
rect 57232 0 57288 400
rect 58576 0 58632 400
rect 59920 0 59976 400
rect 61264 0 61320 400
rect 62608 0 62664 400
rect 63952 0 64008 400
rect 65296 0 65352 400
rect 66640 0 66696 400
rect 67984 0 68040 400
rect 69328 0 69384 400
rect 70672 0 70728 400
rect 72016 0 72072 400
rect 73360 0 73416 400
rect 74704 0 74760 400
rect 76048 0 76104 400
rect 77392 0 77448 400
rect 78736 0 78792 400
rect 80080 0 80136 400
rect 81424 0 81480 400
rect 82768 0 82824 400
rect 84112 0 84168 400
rect 85456 0 85512 400
rect 86800 0 86856 400
rect 88144 0 88200 400
rect 89488 0 89544 400
rect 90832 0 90888 400
rect 92176 0 92232 400
rect 93520 0 93576 400
rect 94864 0 94920 400
rect 96208 0 96264 400
rect 97552 0 97608 400
rect 98896 0 98952 400
rect 100240 0 100296 400
rect 101584 0 101640 400
rect 102928 0 102984 400
rect 104272 0 104328 400
rect 105616 0 105672 400
rect 106960 0 107016 400
rect 108304 0 108360 400
rect 109648 0 109704 400
rect 110992 0 111048 400
rect 112336 0 112392 400
rect 113680 0 113736 400
rect 115024 0 115080 400
rect 116368 0 116424 400
rect 117712 0 117768 400
rect 119056 0 119112 400
rect 120400 0 120456 400
rect 121744 0 121800 400
rect 123088 0 123144 400
rect 124432 0 124488 400
rect 125776 0 125832 400
rect 127120 0 127176 400
rect 128464 0 128520 400
rect 129808 0 129864 400
rect 131152 0 131208 400
rect 132496 0 132552 400
rect 133840 0 133896 400
rect 135184 0 135240 400
rect 136528 0 136584 400
rect 137872 0 137928 400
rect 139216 0 139272 400
rect 140560 0 140616 400
rect 141904 0 141960 400
rect 143248 0 143304 400
rect 144592 0 144648 400
rect 145936 0 145992 400
rect 147280 0 147336 400
rect 148624 0 148680 400
rect 149968 0 150024 400
rect 151312 0 151368 400
rect 152656 0 152712 400
rect 154000 0 154056 400
rect 155344 0 155400 400
rect 156688 0 156744 400
rect 158032 0 158088 400
rect 159376 0 159432 400
rect 160720 0 160776 400
rect 162064 0 162120 400
rect 163408 0 163464 400
rect 164752 0 164808 400
rect 166096 0 166152 400
rect 167440 0 167496 400
rect 168784 0 168840 400
rect 170128 0 170184 400
rect 171472 0 171528 400
rect 172816 0 172872 400
rect 174160 0 174216 400
rect 175504 0 175560 400
rect 176848 0 176904 400
rect 178192 0 178248 400
rect 179536 0 179592 400
rect 180880 0 180936 400
rect 182224 0 182280 400
rect 183568 0 183624 400
rect 184912 0 184968 400
rect 186256 0 186312 400
rect 187600 0 187656 400
rect 188944 0 189000 400
rect 190288 0 190344 400
rect 191632 0 191688 400
rect 192976 0 193032 400
rect 194320 0 194376 400
rect 195664 0 195720 400
rect 197008 0 197064 400
rect 198352 0 198408 400
rect 199696 0 199752 400
rect 201040 0 201096 400
rect 202384 0 202440 400
rect 203728 0 203784 400
rect 205072 0 205128 400
rect 206416 0 206472 400
rect 207760 0 207816 400
rect 209104 0 209160 400
rect 210448 0 210504 400
rect 211792 0 211848 400
rect 213136 0 213192 400
rect 214480 0 214536 400
rect 215824 0 215880 400
rect 217168 0 217224 400
rect 218512 0 218568 400
rect 219856 0 219912 400
rect 221200 0 221256 400
rect 222544 0 222600 400
rect 223888 0 223944 400
rect 225232 0 225288 400
rect 226576 0 226632 400
rect 227920 0 227976 400
rect 229264 0 229320 400
rect 230608 0 230664 400
rect 231952 0 232008 400
rect 233296 0 233352 400
rect 234640 0 234696 400
rect 235984 0 236040 400
rect 237328 0 237384 400
rect 238672 0 238728 400
rect 240016 0 240072 400
rect 241360 0 241416 400
rect 242704 0 242760 400
rect 244048 0 244104 400
rect 245392 0 245448 400
rect 246736 0 246792 400
rect 248080 0 248136 400
rect 249424 0 249480 400
rect 250768 0 250824 400
rect 252112 0 252168 400
rect 253456 0 253512 400
rect 254800 0 254856 400
rect 256144 0 256200 400
rect 257488 0 257544 400
rect 258832 0 258888 400
rect 260176 0 260232 400
rect 261520 0 261576 400
rect 262864 0 262920 400
rect 264208 0 264264 400
rect 265552 0 265608 400
rect 266896 0 266952 400
rect 268240 0 268296 400
rect 269584 0 269640 400
<< obsm2 >>
rect 2238 430 278850 174067
rect 2238 400 10162 430
rect 10278 400 11506 430
rect 11622 400 12850 430
rect 12966 400 14194 430
rect 14310 400 15538 430
rect 15654 400 16882 430
rect 16998 400 18226 430
rect 18342 400 19570 430
rect 19686 400 20914 430
rect 21030 400 22258 430
rect 22374 400 23602 430
rect 23718 400 24946 430
rect 25062 400 26290 430
rect 26406 400 27634 430
rect 27750 400 28978 430
rect 29094 400 30322 430
rect 30438 400 31666 430
rect 31782 400 33010 430
rect 33126 400 34354 430
rect 34470 400 35698 430
rect 35814 400 37042 430
rect 37158 400 38386 430
rect 38502 400 39730 430
rect 39846 400 41074 430
rect 41190 400 42418 430
rect 42534 400 43762 430
rect 43878 400 45106 430
rect 45222 400 46450 430
rect 46566 400 47794 430
rect 47910 400 49138 430
rect 49254 400 50482 430
rect 50598 400 51826 430
rect 51942 400 53170 430
rect 53286 400 54514 430
rect 54630 400 55858 430
rect 55974 400 57202 430
rect 57318 400 58546 430
rect 58662 400 59890 430
rect 60006 400 61234 430
rect 61350 400 62578 430
rect 62694 400 63922 430
rect 64038 400 65266 430
rect 65382 400 66610 430
rect 66726 400 67954 430
rect 68070 400 69298 430
rect 69414 400 70642 430
rect 70758 400 71986 430
rect 72102 400 73330 430
rect 73446 400 74674 430
rect 74790 400 76018 430
rect 76134 400 77362 430
rect 77478 400 78706 430
rect 78822 400 80050 430
rect 80166 400 81394 430
rect 81510 400 82738 430
rect 82854 400 84082 430
rect 84198 400 85426 430
rect 85542 400 86770 430
rect 86886 400 88114 430
rect 88230 400 89458 430
rect 89574 400 90802 430
rect 90918 400 92146 430
rect 92262 400 93490 430
rect 93606 400 94834 430
rect 94950 400 96178 430
rect 96294 400 97522 430
rect 97638 400 98866 430
rect 98982 400 100210 430
rect 100326 400 101554 430
rect 101670 400 102898 430
rect 103014 400 104242 430
rect 104358 400 105586 430
rect 105702 400 106930 430
rect 107046 400 108274 430
rect 108390 400 109618 430
rect 109734 400 110962 430
rect 111078 400 112306 430
rect 112422 400 113650 430
rect 113766 400 114994 430
rect 115110 400 116338 430
rect 116454 400 117682 430
rect 117798 400 119026 430
rect 119142 400 120370 430
rect 120486 400 121714 430
rect 121830 400 123058 430
rect 123174 400 124402 430
rect 124518 400 125746 430
rect 125862 400 127090 430
rect 127206 400 128434 430
rect 128550 400 129778 430
rect 129894 400 131122 430
rect 131238 400 132466 430
rect 132582 400 133810 430
rect 133926 400 135154 430
rect 135270 400 136498 430
rect 136614 400 137842 430
rect 137958 400 139186 430
rect 139302 400 140530 430
rect 140646 400 141874 430
rect 141990 400 143218 430
rect 143334 400 144562 430
rect 144678 400 145906 430
rect 146022 400 147250 430
rect 147366 400 148594 430
rect 148710 400 149938 430
rect 150054 400 151282 430
rect 151398 400 152626 430
rect 152742 400 153970 430
rect 154086 400 155314 430
rect 155430 400 156658 430
rect 156774 400 158002 430
rect 158118 400 159346 430
rect 159462 400 160690 430
rect 160806 400 162034 430
rect 162150 400 163378 430
rect 163494 400 164722 430
rect 164838 400 166066 430
rect 166182 400 167410 430
rect 167526 400 168754 430
rect 168870 400 170098 430
rect 170214 400 171442 430
rect 171558 400 172786 430
rect 172902 400 174130 430
rect 174246 400 175474 430
rect 175590 400 176818 430
rect 176934 400 178162 430
rect 178278 400 179506 430
rect 179622 400 180850 430
rect 180966 400 182194 430
rect 182310 400 183538 430
rect 183654 400 184882 430
rect 184998 400 186226 430
rect 186342 400 187570 430
rect 187686 400 188914 430
rect 189030 400 190258 430
rect 190374 400 191602 430
rect 191718 400 192946 430
rect 193062 400 194290 430
rect 194406 400 195634 430
rect 195750 400 196978 430
rect 197094 400 198322 430
rect 198438 400 199666 430
rect 199782 400 201010 430
rect 201126 400 202354 430
rect 202470 400 203698 430
rect 203814 400 205042 430
rect 205158 400 206386 430
rect 206502 400 207730 430
rect 207846 400 209074 430
rect 209190 400 210418 430
rect 210534 400 211762 430
rect 211878 400 213106 430
rect 213222 400 214450 430
rect 214566 400 215794 430
rect 215910 400 217138 430
rect 217254 400 218482 430
rect 218598 400 219826 430
rect 219942 400 221170 430
rect 221286 400 222514 430
rect 222630 400 223858 430
rect 223974 400 225202 430
rect 225318 400 226546 430
rect 226662 400 227890 430
rect 228006 400 229234 430
rect 229350 400 230578 430
rect 230694 400 231922 430
rect 232038 400 233266 430
rect 233382 400 234610 430
rect 234726 400 235954 430
rect 236070 400 237298 430
rect 237414 400 238642 430
rect 238758 400 239986 430
rect 240102 400 241330 430
rect 241446 400 242674 430
rect 242790 400 244018 430
rect 244134 400 245362 430
rect 245478 400 246706 430
rect 246822 400 248050 430
rect 248166 400 249394 430
rect 249510 400 250738 430
rect 250854 400 252082 430
rect 252198 400 253426 430
rect 253542 400 254770 430
rect 254886 400 256114 430
rect 256230 400 257458 430
rect 257574 400 258802 430
rect 258918 400 260146 430
rect 260262 400 261490 430
rect 261606 400 262834 430
rect 262950 400 264178 430
rect 264294 400 265522 430
rect 265638 400 266866 430
rect 266982 400 268210 430
rect 268326 400 269554 430
rect 269670 400 278850 430
<< obsm3 >>
rect 2233 1554 278855 174062
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< labels >>
rlabel metal2 s 12880 0 12936 400 6 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 53200 0 53256 400 6 la_data_in[10]
port 2 nsew signal input
rlabel metal2 s 57232 0 57288 400 6 la_data_in[11]
port 3 nsew signal input
rlabel metal2 s 61264 0 61320 400 6 la_data_in[12]
port 4 nsew signal input
rlabel metal2 s 65296 0 65352 400 6 la_data_in[13]
port 5 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 la_data_in[14]
port 6 nsew signal input
rlabel metal2 s 73360 0 73416 400 6 la_data_in[15]
port 7 nsew signal input
rlabel metal2 s 77392 0 77448 400 6 la_data_in[16]
port 8 nsew signal input
rlabel metal2 s 81424 0 81480 400 6 la_data_in[17]
port 9 nsew signal input
rlabel metal2 s 85456 0 85512 400 6 la_data_in[18]
port 10 nsew signal input
rlabel metal2 s 89488 0 89544 400 6 la_data_in[19]
port 11 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 la_data_in[1]
port 12 nsew signal input
rlabel metal2 s 93520 0 93576 400 6 la_data_in[20]
port 13 nsew signal input
rlabel metal2 s 97552 0 97608 400 6 la_data_in[21]
port 14 nsew signal input
rlabel metal2 s 101584 0 101640 400 6 la_data_in[22]
port 15 nsew signal input
rlabel metal2 s 105616 0 105672 400 6 la_data_in[23]
port 16 nsew signal input
rlabel metal2 s 109648 0 109704 400 6 la_data_in[24]
port 17 nsew signal input
rlabel metal2 s 113680 0 113736 400 6 la_data_in[25]
port 18 nsew signal input
rlabel metal2 s 117712 0 117768 400 6 la_data_in[26]
port 19 nsew signal input
rlabel metal2 s 121744 0 121800 400 6 la_data_in[27]
port 20 nsew signal input
rlabel metal2 s 125776 0 125832 400 6 la_data_in[28]
port 21 nsew signal input
rlabel metal2 s 129808 0 129864 400 6 la_data_in[29]
port 22 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 la_data_in[2]
port 23 nsew signal input
rlabel metal2 s 133840 0 133896 400 6 la_data_in[30]
port 24 nsew signal input
rlabel metal2 s 137872 0 137928 400 6 la_data_in[31]
port 25 nsew signal input
rlabel metal2 s 141904 0 141960 400 6 la_data_in[32]
port 26 nsew signal input
rlabel metal2 s 145936 0 145992 400 6 la_data_in[33]
port 27 nsew signal input
rlabel metal2 s 149968 0 150024 400 6 la_data_in[34]
port 28 nsew signal input
rlabel metal2 s 154000 0 154056 400 6 la_data_in[35]
port 29 nsew signal input
rlabel metal2 s 158032 0 158088 400 6 la_data_in[36]
port 30 nsew signal input
rlabel metal2 s 162064 0 162120 400 6 la_data_in[37]
port 31 nsew signal input
rlabel metal2 s 166096 0 166152 400 6 la_data_in[38]
port 32 nsew signal input
rlabel metal2 s 170128 0 170184 400 6 la_data_in[39]
port 33 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 la_data_in[3]
port 34 nsew signal input
rlabel metal2 s 174160 0 174216 400 6 la_data_in[40]
port 35 nsew signal input
rlabel metal2 s 178192 0 178248 400 6 la_data_in[41]
port 36 nsew signal input
rlabel metal2 s 182224 0 182280 400 6 la_data_in[42]
port 37 nsew signal input
rlabel metal2 s 186256 0 186312 400 6 la_data_in[43]
port 38 nsew signal input
rlabel metal2 s 190288 0 190344 400 6 la_data_in[44]
port 39 nsew signal input
rlabel metal2 s 194320 0 194376 400 6 la_data_in[45]
port 40 nsew signal input
rlabel metal2 s 198352 0 198408 400 6 la_data_in[46]
port 41 nsew signal input
rlabel metal2 s 202384 0 202440 400 6 la_data_in[47]
port 42 nsew signal input
rlabel metal2 s 206416 0 206472 400 6 la_data_in[48]
port 43 nsew signal input
rlabel metal2 s 210448 0 210504 400 6 la_data_in[49]
port 44 nsew signal input
rlabel metal2 s 29008 0 29064 400 6 la_data_in[4]
port 45 nsew signal input
rlabel metal2 s 214480 0 214536 400 6 la_data_in[50]
port 46 nsew signal input
rlabel metal2 s 218512 0 218568 400 6 la_data_in[51]
port 47 nsew signal input
rlabel metal2 s 222544 0 222600 400 6 la_data_in[52]
port 48 nsew signal input
rlabel metal2 s 226576 0 226632 400 6 la_data_in[53]
port 49 nsew signal input
rlabel metal2 s 230608 0 230664 400 6 la_data_in[54]
port 50 nsew signal input
rlabel metal2 s 234640 0 234696 400 6 la_data_in[55]
port 51 nsew signal input
rlabel metal2 s 238672 0 238728 400 6 la_data_in[56]
port 52 nsew signal input
rlabel metal2 s 242704 0 242760 400 6 la_data_in[57]
port 53 nsew signal input
rlabel metal2 s 246736 0 246792 400 6 la_data_in[58]
port 54 nsew signal input
rlabel metal2 s 250768 0 250824 400 6 la_data_in[59]
port 55 nsew signal input
rlabel metal2 s 33040 0 33096 400 6 la_data_in[5]
port 56 nsew signal input
rlabel metal2 s 254800 0 254856 400 6 la_data_in[60]
port 57 nsew signal input
rlabel metal2 s 258832 0 258888 400 6 la_data_in[61]
port 58 nsew signal input
rlabel metal2 s 262864 0 262920 400 6 la_data_in[62]
port 59 nsew signal input
rlabel metal2 s 266896 0 266952 400 6 la_data_in[63]
port 60 nsew signal input
rlabel metal2 s 37072 0 37128 400 6 la_data_in[6]
port 61 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 la_data_in[7]
port 62 nsew signal input
rlabel metal2 s 45136 0 45192 400 6 la_data_in[8]
port 63 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 la_data_in[9]
port 64 nsew signal input
rlabel metal2 s 14224 0 14280 400 6 la_data_out[0]
port 65 nsew signal output
rlabel metal2 s 54544 0 54600 400 6 la_data_out[10]
port 66 nsew signal output
rlabel metal2 s 58576 0 58632 400 6 la_data_out[11]
port 67 nsew signal output
rlabel metal2 s 62608 0 62664 400 6 la_data_out[12]
port 68 nsew signal output
rlabel metal2 s 66640 0 66696 400 6 la_data_out[13]
port 69 nsew signal output
rlabel metal2 s 70672 0 70728 400 6 la_data_out[14]
port 70 nsew signal output
rlabel metal2 s 74704 0 74760 400 6 la_data_out[15]
port 71 nsew signal output
rlabel metal2 s 78736 0 78792 400 6 la_data_out[16]
port 72 nsew signal output
rlabel metal2 s 82768 0 82824 400 6 la_data_out[17]
port 73 nsew signal output
rlabel metal2 s 86800 0 86856 400 6 la_data_out[18]
port 74 nsew signal output
rlabel metal2 s 90832 0 90888 400 6 la_data_out[19]
port 75 nsew signal output
rlabel metal2 s 18256 0 18312 400 6 la_data_out[1]
port 76 nsew signal output
rlabel metal2 s 94864 0 94920 400 6 la_data_out[20]
port 77 nsew signal output
rlabel metal2 s 98896 0 98952 400 6 la_data_out[21]
port 78 nsew signal output
rlabel metal2 s 102928 0 102984 400 6 la_data_out[22]
port 79 nsew signal output
rlabel metal2 s 106960 0 107016 400 6 la_data_out[23]
port 80 nsew signal output
rlabel metal2 s 110992 0 111048 400 6 la_data_out[24]
port 81 nsew signal output
rlabel metal2 s 115024 0 115080 400 6 la_data_out[25]
port 82 nsew signal output
rlabel metal2 s 119056 0 119112 400 6 la_data_out[26]
port 83 nsew signal output
rlabel metal2 s 123088 0 123144 400 6 la_data_out[27]
port 84 nsew signal output
rlabel metal2 s 127120 0 127176 400 6 la_data_out[28]
port 85 nsew signal output
rlabel metal2 s 131152 0 131208 400 6 la_data_out[29]
port 86 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 la_data_out[2]
port 87 nsew signal output
rlabel metal2 s 135184 0 135240 400 6 la_data_out[30]
port 88 nsew signal output
rlabel metal2 s 139216 0 139272 400 6 la_data_out[31]
port 89 nsew signal output
rlabel metal2 s 143248 0 143304 400 6 la_data_out[32]
port 90 nsew signal output
rlabel metal2 s 147280 0 147336 400 6 la_data_out[33]
port 91 nsew signal output
rlabel metal2 s 151312 0 151368 400 6 la_data_out[34]
port 92 nsew signal output
rlabel metal2 s 155344 0 155400 400 6 la_data_out[35]
port 93 nsew signal output
rlabel metal2 s 159376 0 159432 400 6 la_data_out[36]
port 94 nsew signal output
rlabel metal2 s 163408 0 163464 400 6 la_data_out[37]
port 95 nsew signal output
rlabel metal2 s 167440 0 167496 400 6 la_data_out[38]
port 96 nsew signal output
rlabel metal2 s 171472 0 171528 400 6 la_data_out[39]
port 97 nsew signal output
rlabel metal2 s 26320 0 26376 400 6 la_data_out[3]
port 98 nsew signal output
rlabel metal2 s 175504 0 175560 400 6 la_data_out[40]
port 99 nsew signal output
rlabel metal2 s 179536 0 179592 400 6 la_data_out[41]
port 100 nsew signal output
rlabel metal2 s 183568 0 183624 400 6 la_data_out[42]
port 101 nsew signal output
rlabel metal2 s 187600 0 187656 400 6 la_data_out[43]
port 102 nsew signal output
rlabel metal2 s 191632 0 191688 400 6 la_data_out[44]
port 103 nsew signal output
rlabel metal2 s 195664 0 195720 400 6 la_data_out[45]
port 104 nsew signal output
rlabel metal2 s 199696 0 199752 400 6 la_data_out[46]
port 105 nsew signal output
rlabel metal2 s 203728 0 203784 400 6 la_data_out[47]
port 106 nsew signal output
rlabel metal2 s 207760 0 207816 400 6 la_data_out[48]
port 107 nsew signal output
rlabel metal2 s 211792 0 211848 400 6 la_data_out[49]
port 108 nsew signal output
rlabel metal2 s 30352 0 30408 400 6 la_data_out[4]
port 109 nsew signal output
rlabel metal2 s 215824 0 215880 400 6 la_data_out[50]
port 110 nsew signal output
rlabel metal2 s 219856 0 219912 400 6 la_data_out[51]
port 111 nsew signal output
rlabel metal2 s 223888 0 223944 400 6 la_data_out[52]
port 112 nsew signal output
rlabel metal2 s 227920 0 227976 400 6 la_data_out[53]
port 113 nsew signal output
rlabel metal2 s 231952 0 232008 400 6 la_data_out[54]
port 114 nsew signal output
rlabel metal2 s 235984 0 236040 400 6 la_data_out[55]
port 115 nsew signal output
rlabel metal2 s 240016 0 240072 400 6 la_data_out[56]
port 116 nsew signal output
rlabel metal2 s 244048 0 244104 400 6 la_data_out[57]
port 117 nsew signal output
rlabel metal2 s 248080 0 248136 400 6 la_data_out[58]
port 118 nsew signal output
rlabel metal2 s 252112 0 252168 400 6 la_data_out[59]
port 119 nsew signal output
rlabel metal2 s 34384 0 34440 400 6 la_data_out[5]
port 120 nsew signal output
rlabel metal2 s 256144 0 256200 400 6 la_data_out[60]
port 121 nsew signal output
rlabel metal2 s 260176 0 260232 400 6 la_data_out[61]
port 122 nsew signal output
rlabel metal2 s 264208 0 264264 400 6 la_data_out[62]
port 123 nsew signal output
rlabel metal2 s 268240 0 268296 400 6 la_data_out[63]
port 124 nsew signal output
rlabel metal2 s 38416 0 38472 400 6 la_data_out[6]
port 125 nsew signal output
rlabel metal2 s 42448 0 42504 400 6 la_data_out[7]
port 126 nsew signal output
rlabel metal2 s 46480 0 46536 400 6 la_data_out[8]
port 127 nsew signal output
rlabel metal2 s 50512 0 50568 400 6 la_data_out[9]
port 128 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 la_oenb[0]
port 129 nsew signal input
rlabel metal2 s 55888 0 55944 400 6 la_oenb[10]
port 130 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 la_oenb[11]
port 131 nsew signal input
rlabel metal2 s 63952 0 64008 400 6 la_oenb[12]
port 132 nsew signal input
rlabel metal2 s 67984 0 68040 400 6 la_oenb[13]
port 133 nsew signal input
rlabel metal2 s 72016 0 72072 400 6 la_oenb[14]
port 134 nsew signal input
rlabel metal2 s 76048 0 76104 400 6 la_oenb[15]
port 135 nsew signal input
rlabel metal2 s 80080 0 80136 400 6 la_oenb[16]
port 136 nsew signal input
rlabel metal2 s 84112 0 84168 400 6 la_oenb[17]
port 137 nsew signal input
rlabel metal2 s 88144 0 88200 400 6 la_oenb[18]
port 138 nsew signal input
rlabel metal2 s 92176 0 92232 400 6 la_oenb[19]
port 139 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 la_oenb[1]
port 140 nsew signal input
rlabel metal2 s 96208 0 96264 400 6 la_oenb[20]
port 141 nsew signal input
rlabel metal2 s 100240 0 100296 400 6 la_oenb[21]
port 142 nsew signal input
rlabel metal2 s 104272 0 104328 400 6 la_oenb[22]
port 143 nsew signal input
rlabel metal2 s 108304 0 108360 400 6 la_oenb[23]
port 144 nsew signal input
rlabel metal2 s 112336 0 112392 400 6 la_oenb[24]
port 145 nsew signal input
rlabel metal2 s 116368 0 116424 400 6 la_oenb[25]
port 146 nsew signal input
rlabel metal2 s 120400 0 120456 400 6 la_oenb[26]
port 147 nsew signal input
rlabel metal2 s 124432 0 124488 400 6 la_oenb[27]
port 148 nsew signal input
rlabel metal2 s 128464 0 128520 400 6 la_oenb[28]
port 149 nsew signal input
rlabel metal2 s 132496 0 132552 400 6 la_oenb[29]
port 150 nsew signal input
rlabel metal2 s 23632 0 23688 400 6 la_oenb[2]
port 151 nsew signal input
rlabel metal2 s 136528 0 136584 400 6 la_oenb[30]
port 152 nsew signal input
rlabel metal2 s 140560 0 140616 400 6 la_oenb[31]
port 153 nsew signal input
rlabel metal2 s 144592 0 144648 400 6 la_oenb[32]
port 154 nsew signal input
rlabel metal2 s 148624 0 148680 400 6 la_oenb[33]
port 155 nsew signal input
rlabel metal2 s 152656 0 152712 400 6 la_oenb[34]
port 156 nsew signal input
rlabel metal2 s 156688 0 156744 400 6 la_oenb[35]
port 157 nsew signal input
rlabel metal2 s 160720 0 160776 400 6 la_oenb[36]
port 158 nsew signal input
rlabel metal2 s 164752 0 164808 400 6 la_oenb[37]
port 159 nsew signal input
rlabel metal2 s 168784 0 168840 400 6 la_oenb[38]
port 160 nsew signal input
rlabel metal2 s 172816 0 172872 400 6 la_oenb[39]
port 161 nsew signal input
rlabel metal2 s 27664 0 27720 400 6 la_oenb[3]
port 162 nsew signal input
rlabel metal2 s 176848 0 176904 400 6 la_oenb[40]
port 163 nsew signal input
rlabel metal2 s 180880 0 180936 400 6 la_oenb[41]
port 164 nsew signal input
rlabel metal2 s 184912 0 184968 400 6 la_oenb[42]
port 165 nsew signal input
rlabel metal2 s 188944 0 189000 400 6 la_oenb[43]
port 166 nsew signal input
rlabel metal2 s 192976 0 193032 400 6 la_oenb[44]
port 167 nsew signal input
rlabel metal2 s 197008 0 197064 400 6 la_oenb[45]
port 168 nsew signal input
rlabel metal2 s 201040 0 201096 400 6 la_oenb[46]
port 169 nsew signal input
rlabel metal2 s 205072 0 205128 400 6 la_oenb[47]
port 170 nsew signal input
rlabel metal2 s 209104 0 209160 400 6 la_oenb[48]
port 171 nsew signal input
rlabel metal2 s 213136 0 213192 400 6 la_oenb[49]
port 172 nsew signal input
rlabel metal2 s 31696 0 31752 400 6 la_oenb[4]
port 173 nsew signal input
rlabel metal2 s 217168 0 217224 400 6 la_oenb[50]
port 174 nsew signal input
rlabel metal2 s 221200 0 221256 400 6 la_oenb[51]
port 175 nsew signal input
rlabel metal2 s 225232 0 225288 400 6 la_oenb[52]
port 176 nsew signal input
rlabel metal2 s 229264 0 229320 400 6 la_oenb[53]
port 177 nsew signal input
rlabel metal2 s 233296 0 233352 400 6 la_oenb[54]
port 178 nsew signal input
rlabel metal2 s 237328 0 237384 400 6 la_oenb[55]
port 179 nsew signal input
rlabel metal2 s 241360 0 241416 400 6 la_oenb[56]
port 180 nsew signal input
rlabel metal2 s 245392 0 245448 400 6 la_oenb[57]
port 181 nsew signal input
rlabel metal2 s 249424 0 249480 400 6 la_oenb[58]
port 182 nsew signal input
rlabel metal2 s 253456 0 253512 400 6 la_oenb[59]
port 183 nsew signal input
rlabel metal2 s 35728 0 35784 400 6 la_oenb[5]
port 184 nsew signal input
rlabel metal2 s 257488 0 257544 400 6 la_oenb[60]
port 185 nsew signal input
rlabel metal2 s 261520 0 261576 400 6 la_oenb[61]
port 186 nsew signal input
rlabel metal2 s 265552 0 265608 400 6 la_oenb[62]
port 187 nsew signal input
rlabel metal2 s 269584 0 269640 400 6 la_oenb[63]
port 188 nsew signal input
rlabel metal2 s 39760 0 39816 400 6 la_oenb[6]
port 189 nsew signal input
rlabel metal2 s 43792 0 43848 400 6 la_oenb[7]
port 190 nsew signal input
rlabel metal2 s 47824 0 47880 400 6 la_oenb[8]
port 191 nsew signal input
rlabel metal2 s 51856 0 51912 400 6 la_oenb[9]
port 192 nsew signal input
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 193 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 194 nsew ground bidirectional
rlabel metal2 s 10192 0 10248 400 6 wb_clk_i
port 195 nsew signal input
rlabel metal2 s 11536 0 11592 400 6 wb_rst_i
port 196 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14916238
string GDS_FILE /home/hiepdm/hello/openlane/user_proj_example/runs/23_12_10_08_16/results/signoff/user_proj_example.magic.gds
string GDS_START 49130
<< end >>

