VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 572.320 0.000 572.880 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 612.640 0.000 613.200 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 652.960 0.000 653.520 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 0.000 693.840 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 733.600 0.000 734.160 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 773.920 0.000 774.480 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 814.240 0.000 814.800 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 854.560 0.000 855.120 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 894.880 0.000 895.440 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 935.200 0.000 935.760 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 975.520 0.000 976.080 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1015.840 0.000 1016.400 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.160 0.000 1056.720 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1096.480 0.000 1097.040 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1136.800 0.000 1137.360 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1177.120 0.000 1177.680 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1217.440 0.000 1218.000 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1257.760 0.000 1258.320 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1298.080 0.000 1298.640 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1338.400 0.000 1338.960 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1378.720 0.000 1379.280 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1419.040 0.000 1419.600 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1459.360 0.000 1459.920 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1499.680 0.000 1500.240 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1540.000 0.000 1540.560 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1580.320 0.000 1580.880 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1620.640 0.000 1621.200 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1660.960 0.000 1661.520 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1701.280 0.000 1701.840 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1741.600 0.000 1742.160 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1781.920 0.000 1782.480 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1822.240 0.000 1822.800 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1862.560 0.000 1863.120 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1902.880 0.000 1903.440 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1943.200 0.000 1943.760 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1983.520 0.000 1984.080 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2023.840 0.000 2024.400 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2064.160 0.000 2064.720 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2104.480 0.000 2105.040 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2144.800 0.000 2145.360 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2185.120 0.000 2185.680 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2225.440 0.000 2226.000 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2265.760 0.000 2266.320 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2306.080 0.000 2306.640 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2346.400 0.000 2346.960 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2386.720 0.000 2387.280 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2427.040 0.000 2427.600 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2467.360 0.000 2467.920 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2507.680 0.000 2508.240 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 0.000 330.960 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2548.000 0.000 2548.560 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2588.320 0.000 2588.880 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2628.640 0.000 2629.200 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2668.960 0.000 2669.520 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 0.000 371.280 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 0.000 411.600 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 0.000 451.920 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 0.000 492.240 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 545.440 0.000 546.000 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 585.760 0.000 586.320 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 0.000 626.640 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 666.400 0.000 666.960 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 0.000 707.280 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 747.040 0.000 747.600 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 787.360 0.000 787.920 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 0.000 828.240 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 868.000 0.000 868.560 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 908.320 0.000 908.880 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 948.640 0.000 949.200 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 988.960 0.000 989.520 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1029.280 0.000 1029.840 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1069.600 0.000 1070.160 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1109.920 0.000 1110.480 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1150.240 0.000 1150.800 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1190.560 0.000 1191.120 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1230.880 0.000 1231.440 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1271.200 0.000 1271.760 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1311.520 0.000 1312.080 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1351.840 0.000 1352.400 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1392.160 0.000 1392.720 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1432.480 0.000 1433.040 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1472.800 0.000 1473.360 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1513.120 0.000 1513.680 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1553.440 0.000 1554.000 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1593.760 0.000 1594.320 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1634.080 0.000 1634.640 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1674.400 0.000 1674.960 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1714.720 0.000 1715.280 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1755.040 0.000 1755.600 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1795.360 0.000 1795.920 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1835.680 0.000 1836.240 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1876.000 0.000 1876.560 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1916.320 0.000 1916.880 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1956.640 0.000 1957.200 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1996.960 0.000 1997.520 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2037.280 0.000 2037.840 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2077.600 0.000 2078.160 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2117.920 0.000 2118.480 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 0.000 304.080 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2158.240 0.000 2158.800 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2198.560 0.000 2199.120 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2238.880 0.000 2239.440 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2279.200 0.000 2279.760 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2319.520 0.000 2320.080 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2359.840 0.000 2360.400 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2400.160 0.000 2400.720 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2440.480 0.000 2441.040 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2480.800 0.000 2481.360 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2521.120 0.000 2521.680 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 0.000 344.400 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2561.440 0.000 2562.000 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2601.760 0.000 2602.320 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2642.080 0.000 2642.640 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2682.400 0.000 2682.960 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 384.160 0.000 384.720 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 0.000 465.360 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 0.000 505.680 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 0.000 559.440 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 0.000 599.760 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 0.000 640.080 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 679.840 0.000 680.400 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 0.000 720.720 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 0.000 761.040 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 800.800 0.000 801.360 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 0.000 841.680 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 881.440 0.000 882.000 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 921.760 0.000 922.320 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 0.000 962.640 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1002.400 0.000 1002.960 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1042.720 0.000 1043.280 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1083.040 0.000 1083.600 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1123.360 0.000 1123.920 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1163.680 0.000 1164.240 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1204.000 0.000 1204.560 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1244.320 0.000 1244.880 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1284.640 0.000 1285.200 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1324.960 0.000 1325.520 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 0.000 236.880 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1365.280 0.000 1365.840 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1405.600 0.000 1406.160 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1445.920 0.000 1446.480 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1486.240 0.000 1486.800 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1526.560 0.000 1527.120 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1566.880 0.000 1567.440 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1607.200 0.000 1607.760 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1647.520 0.000 1648.080 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1687.840 0.000 1688.400 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1728.160 0.000 1728.720 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1768.480 0.000 1769.040 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1808.800 0.000 1809.360 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1849.120 0.000 1849.680 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1889.440 0.000 1890.000 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1929.760 0.000 1930.320 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1970.080 0.000 1970.640 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2010.400 0.000 2010.960 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2050.720 0.000 2051.280 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2091.040 0.000 2091.600 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2131.360 0.000 2131.920 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 0.000 317.520 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2171.680 0.000 2172.240 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2212.000 0.000 2212.560 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2252.320 0.000 2252.880 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2292.640 0.000 2293.200 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2332.960 0.000 2333.520 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2373.280 0.000 2373.840 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2413.600 0.000 2414.160 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2453.920 0.000 2454.480 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2494.240 0.000 2494.800 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2534.560 0.000 2535.120 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2574.880 0.000 2575.440 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2615.200 0.000 2615.760 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2655.520 0.000 2656.080 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2695.840 0.000 2696.400 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 0.000 398.160 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 0.000 438.480 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 0.000 478.800 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 0.000 519.120 4.000 ;
    END
  END la_oenb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1740.780 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1740.780 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER Pwell ;
        RECT 6.290 1738.720 2793.710 1740.910 ;
      LAYER Nwell ;
        RECT 6.290 1734.400 2793.710 1738.720 ;
      LAYER Pwell ;
        RECT 6.290 1730.880 2793.710 1734.400 ;
      LAYER Nwell ;
        RECT 6.290 1726.560 2793.710 1730.880 ;
      LAYER Pwell ;
        RECT 6.290 1723.040 2793.710 1726.560 ;
      LAYER Nwell ;
        RECT 6.290 1718.720 2793.710 1723.040 ;
      LAYER Pwell ;
        RECT 6.290 1715.200 2793.710 1718.720 ;
      LAYER Nwell ;
        RECT 6.290 1710.880 2793.710 1715.200 ;
      LAYER Pwell ;
        RECT 6.290 1707.360 2793.710 1710.880 ;
      LAYER Nwell ;
        RECT 6.290 1703.040 2793.710 1707.360 ;
      LAYER Pwell ;
        RECT 6.290 1699.520 2793.710 1703.040 ;
      LAYER Nwell ;
        RECT 6.290 1695.200 2793.710 1699.520 ;
      LAYER Pwell ;
        RECT 6.290 1691.680 2793.710 1695.200 ;
      LAYER Nwell ;
        RECT 6.290 1687.360 2793.710 1691.680 ;
      LAYER Pwell ;
        RECT 6.290 1683.840 2793.710 1687.360 ;
      LAYER Nwell ;
        RECT 6.290 1679.520 2793.710 1683.840 ;
      LAYER Pwell ;
        RECT 6.290 1676.000 2793.710 1679.520 ;
      LAYER Nwell ;
        RECT 6.290 1671.680 2793.710 1676.000 ;
      LAYER Pwell ;
        RECT 6.290 1668.160 2793.710 1671.680 ;
      LAYER Nwell ;
        RECT 6.290 1663.840 2793.710 1668.160 ;
      LAYER Pwell ;
        RECT 6.290 1660.320 2793.710 1663.840 ;
      LAYER Nwell ;
        RECT 6.290 1656.000 2793.710 1660.320 ;
      LAYER Pwell ;
        RECT 6.290 1652.480 2793.710 1656.000 ;
      LAYER Nwell ;
        RECT 6.290 1648.160 2793.710 1652.480 ;
      LAYER Pwell ;
        RECT 6.290 1644.640 2793.710 1648.160 ;
      LAYER Nwell ;
        RECT 6.290 1640.320 2793.710 1644.640 ;
      LAYER Pwell ;
        RECT 6.290 1636.800 2793.710 1640.320 ;
      LAYER Nwell ;
        RECT 6.290 1632.480 2793.710 1636.800 ;
      LAYER Pwell ;
        RECT 6.290 1628.960 2793.710 1632.480 ;
      LAYER Nwell ;
        RECT 6.290 1624.640 2793.710 1628.960 ;
      LAYER Pwell ;
        RECT 6.290 1621.120 2793.710 1624.640 ;
      LAYER Nwell ;
        RECT 6.290 1616.800 2793.710 1621.120 ;
      LAYER Pwell ;
        RECT 6.290 1613.280 2793.710 1616.800 ;
      LAYER Nwell ;
        RECT 6.290 1608.960 2793.710 1613.280 ;
      LAYER Pwell ;
        RECT 6.290 1605.440 2793.710 1608.960 ;
      LAYER Nwell ;
        RECT 6.290 1601.120 2793.710 1605.440 ;
      LAYER Pwell ;
        RECT 6.290 1597.600 2793.710 1601.120 ;
      LAYER Nwell ;
        RECT 6.290 1593.280 2793.710 1597.600 ;
      LAYER Pwell ;
        RECT 6.290 1589.760 2793.710 1593.280 ;
      LAYER Nwell ;
        RECT 6.290 1585.440 2793.710 1589.760 ;
      LAYER Pwell ;
        RECT 6.290 1581.920 2793.710 1585.440 ;
      LAYER Nwell ;
        RECT 6.290 1577.600 2793.710 1581.920 ;
      LAYER Pwell ;
        RECT 6.290 1574.080 2793.710 1577.600 ;
      LAYER Nwell ;
        RECT 6.290 1569.760 2793.710 1574.080 ;
      LAYER Pwell ;
        RECT 6.290 1566.240 2793.710 1569.760 ;
      LAYER Nwell ;
        RECT 6.290 1561.920 2793.710 1566.240 ;
      LAYER Pwell ;
        RECT 6.290 1558.400 2793.710 1561.920 ;
      LAYER Nwell ;
        RECT 6.290 1554.080 2793.710 1558.400 ;
      LAYER Pwell ;
        RECT 6.290 1550.560 2793.710 1554.080 ;
      LAYER Nwell ;
        RECT 6.290 1546.240 2793.710 1550.560 ;
      LAYER Pwell ;
        RECT 6.290 1542.720 2793.710 1546.240 ;
      LAYER Nwell ;
        RECT 6.290 1538.400 2793.710 1542.720 ;
      LAYER Pwell ;
        RECT 6.290 1534.880 2793.710 1538.400 ;
      LAYER Nwell ;
        RECT 6.290 1530.560 2793.710 1534.880 ;
      LAYER Pwell ;
        RECT 6.290 1527.040 2793.710 1530.560 ;
      LAYER Nwell ;
        RECT 6.290 1522.720 2793.710 1527.040 ;
      LAYER Pwell ;
        RECT 6.290 1519.200 2793.710 1522.720 ;
      LAYER Nwell ;
        RECT 6.290 1514.880 2793.710 1519.200 ;
      LAYER Pwell ;
        RECT 6.290 1511.360 2793.710 1514.880 ;
      LAYER Nwell ;
        RECT 6.290 1507.040 2793.710 1511.360 ;
      LAYER Pwell ;
        RECT 6.290 1503.520 2793.710 1507.040 ;
      LAYER Nwell ;
        RECT 6.290 1499.200 2793.710 1503.520 ;
      LAYER Pwell ;
        RECT 6.290 1495.680 2793.710 1499.200 ;
      LAYER Nwell ;
        RECT 6.290 1491.360 2793.710 1495.680 ;
      LAYER Pwell ;
        RECT 6.290 1487.840 2793.710 1491.360 ;
      LAYER Nwell ;
        RECT 6.290 1483.520 2793.710 1487.840 ;
      LAYER Pwell ;
        RECT 6.290 1480.000 2793.710 1483.520 ;
      LAYER Nwell ;
        RECT 6.290 1475.680 2793.710 1480.000 ;
      LAYER Pwell ;
        RECT 6.290 1472.160 2793.710 1475.680 ;
      LAYER Nwell ;
        RECT 6.290 1467.840 2793.710 1472.160 ;
      LAYER Pwell ;
        RECT 6.290 1464.320 2793.710 1467.840 ;
      LAYER Nwell ;
        RECT 6.290 1460.000 2793.710 1464.320 ;
      LAYER Pwell ;
        RECT 6.290 1456.480 2793.710 1460.000 ;
      LAYER Nwell ;
        RECT 6.290 1452.160 2793.710 1456.480 ;
      LAYER Pwell ;
        RECT 6.290 1448.640 2793.710 1452.160 ;
      LAYER Nwell ;
        RECT 6.290 1444.320 2793.710 1448.640 ;
      LAYER Pwell ;
        RECT 6.290 1440.800 2793.710 1444.320 ;
      LAYER Nwell ;
        RECT 6.290 1436.480 2793.710 1440.800 ;
      LAYER Pwell ;
        RECT 6.290 1432.960 2793.710 1436.480 ;
      LAYER Nwell ;
        RECT 6.290 1428.640 2793.710 1432.960 ;
      LAYER Pwell ;
        RECT 6.290 1425.120 2793.710 1428.640 ;
      LAYER Nwell ;
        RECT 6.290 1420.800 2793.710 1425.120 ;
      LAYER Pwell ;
        RECT 6.290 1417.280 2793.710 1420.800 ;
      LAYER Nwell ;
        RECT 6.290 1412.960 2793.710 1417.280 ;
      LAYER Pwell ;
        RECT 6.290 1409.440 2793.710 1412.960 ;
      LAYER Nwell ;
        RECT 6.290 1405.120 2793.710 1409.440 ;
      LAYER Pwell ;
        RECT 6.290 1401.600 2793.710 1405.120 ;
      LAYER Nwell ;
        RECT 6.290 1397.280 2793.710 1401.600 ;
      LAYER Pwell ;
        RECT 6.290 1393.760 2793.710 1397.280 ;
      LAYER Nwell ;
        RECT 6.290 1389.440 2793.710 1393.760 ;
      LAYER Pwell ;
        RECT 6.290 1385.920 2793.710 1389.440 ;
      LAYER Nwell ;
        RECT 6.290 1381.600 2793.710 1385.920 ;
      LAYER Pwell ;
        RECT 6.290 1378.080 2793.710 1381.600 ;
      LAYER Nwell ;
        RECT 6.290 1373.760 2793.710 1378.080 ;
      LAYER Pwell ;
        RECT 6.290 1370.240 2793.710 1373.760 ;
      LAYER Nwell ;
        RECT 6.290 1365.920 2793.710 1370.240 ;
      LAYER Pwell ;
        RECT 6.290 1362.400 2793.710 1365.920 ;
      LAYER Nwell ;
        RECT 6.290 1358.080 2793.710 1362.400 ;
      LAYER Pwell ;
        RECT 6.290 1354.560 2793.710 1358.080 ;
      LAYER Nwell ;
        RECT 6.290 1350.240 2793.710 1354.560 ;
      LAYER Pwell ;
        RECT 6.290 1346.720 2793.710 1350.240 ;
      LAYER Nwell ;
        RECT 6.290 1342.400 2793.710 1346.720 ;
      LAYER Pwell ;
        RECT 6.290 1338.880 2793.710 1342.400 ;
      LAYER Nwell ;
        RECT 6.290 1334.560 2793.710 1338.880 ;
      LAYER Pwell ;
        RECT 6.290 1331.040 2793.710 1334.560 ;
      LAYER Nwell ;
        RECT 6.290 1326.720 2793.710 1331.040 ;
      LAYER Pwell ;
        RECT 6.290 1323.200 2793.710 1326.720 ;
      LAYER Nwell ;
        RECT 6.290 1318.880 2793.710 1323.200 ;
      LAYER Pwell ;
        RECT 6.290 1315.360 2793.710 1318.880 ;
      LAYER Nwell ;
        RECT 6.290 1311.040 2793.710 1315.360 ;
      LAYER Pwell ;
        RECT 6.290 1307.520 2793.710 1311.040 ;
      LAYER Nwell ;
        RECT 6.290 1303.200 2793.710 1307.520 ;
      LAYER Pwell ;
        RECT 6.290 1299.680 2793.710 1303.200 ;
      LAYER Nwell ;
        RECT 6.290 1295.360 2793.710 1299.680 ;
      LAYER Pwell ;
        RECT 6.290 1291.840 2793.710 1295.360 ;
      LAYER Nwell ;
        RECT 6.290 1287.520 2793.710 1291.840 ;
      LAYER Pwell ;
        RECT 6.290 1284.000 2793.710 1287.520 ;
      LAYER Nwell ;
        RECT 6.290 1279.680 2793.710 1284.000 ;
      LAYER Pwell ;
        RECT 6.290 1276.160 2793.710 1279.680 ;
      LAYER Nwell ;
        RECT 6.290 1271.840 2793.710 1276.160 ;
      LAYER Pwell ;
        RECT 6.290 1268.320 2793.710 1271.840 ;
      LAYER Nwell ;
        RECT 6.290 1264.000 2793.710 1268.320 ;
      LAYER Pwell ;
        RECT 6.290 1260.480 2793.710 1264.000 ;
      LAYER Nwell ;
        RECT 6.290 1256.160 2793.710 1260.480 ;
      LAYER Pwell ;
        RECT 6.290 1252.640 2793.710 1256.160 ;
      LAYER Nwell ;
        RECT 6.290 1248.320 2793.710 1252.640 ;
      LAYER Pwell ;
        RECT 6.290 1244.800 2793.710 1248.320 ;
      LAYER Nwell ;
        RECT 6.290 1240.480 2793.710 1244.800 ;
      LAYER Pwell ;
        RECT 6.290 1236.960 2793.710 1240.480 ;
      LAYER Nwell ;
        RECT 6.290 1232.640 2793.710 1236.960 ;
      LAYER Pwell ;
        RECT 6.290 1229.120 2793.710 1232.640 ;
      LAYER Nwell ;
        RECT 6.290 1224.800 2793.710 1229.120 ;
      LAYER Pwell ;
        RECT 6.290 1221.280 2793.710 1224.800 ;
      LAYER Nwell ;
        RECT 6.290 1216.960 2793.710 1221.280 ;
      LAYER Pwell ;
        RECT 6.290 1213.440 2793.710 1216.960 ;
      LAYER Nwell ;
        RECT 6.290 1209.120 2793.710 1213.440 ;
      LAYER Pwell ;
        RECT 6.290 1205.600 2793.710 1209.120 ;
      LAYER Nwell ;
        RECT 6.290 1201.280 2793.710 1205.600 ;
      LAYER Pwell ;
        RECT 6.290 1197.760 2793.710 1201.280 ;
      LAYER Nwell ;
        RECT 6.290 1193.440 2793.710 1197.760 ;
      LAYER Pwell ;
        RECT 6.290 1189.920 2793.710 1193.440 ;
      LAYER Nwell ;
        RECT 6.290 1185.600 2793.710 1189.920 ;
      LAYER Pwell ;
        RECT 6.290 1182.080 2793.710 1185.600 ;
      LAYER Nwell ;
        RECT 6.290 1177.760 2793.710 1182.080 ;
      LAYER Pwell ;
        RECT 6.290 1174.240 2793.710 1177.760 ;
      LAYER Nwell ;
        RECT 6.290 1169.920 2793.710 1174.240 ;
      LAYER Pwell ;
        RECT 6.290 1166.400 2793.710 1169.920 ;
      LAYER Nwell ;
        RECT 6.290 1162.080 2793.710 1166.400 ;
      LAYER Pwell ;
        RECT 6.290 1158.560 2793.710 1162.080 ;
      LAYER Nwell ;
        RECT 6.290 1154.240 2793.710 1158.560 ;
      LAYER Pwell ;
        RECT 6.290 1150.720 2793.710 1154.240 ;
      LAYER Nwell ;
        RECT 6.290 1146.400 2793.710 1150.720 ;
      LAYER Pwell ;
        RECT 6.290 1142.880 2793.710 1146.400 ;
      LAYER Nwell ;
        RECT 6.290 1138.560 2793.710 1142.880 ;
      LAYER Pwell ;
        RECT 6.290 1135.040 2793.710 1138.560 ;
      LAYER Nwell ;
        RECT 6.290 1130.720 2793.710 1135.040 ;
      LAYER Pwell ;
        RECT 6.290 1127.200 2793.710 1130.720 ;
      LAYER Nwell ;
        RECT 6.290 1122.880 2793.710 1127.200 ;
      LAYER Pwell ;
        RECT 6.290 1119.360 2793.710 1122.880 ;
      LAYER Nwell ;
        RECT 6.290 1115.040 2793.710 1119.360 ;
      LAYER Pwell ;
        RECT 6.290 1111.520 2793.710 1115.040 ;
      LAYER Nwell ;
        RECT 6.290 1107.200 2793.710 1111.520 ;
      LAYER Pwell ;
        RECT 6.290 1103.680 2793.710 1107.200 ;
      LAYER Nwell ;
        RECT 6.290 1099.360 2793.710 1103.680 ;
      LAYER Pwell ;
        RECT 6.290 1095.840 2793.710 1099.360 ;
      LAYER Nwell ;
        RECT 6.290 1091.520 2793.710 1095.840 ;
      LAYER Pwell ;
        RECT 6.290 1088.000 2793.710 1091.520 ;
      LAYER Nwell ;
        RECT 6.290 1083.680 2793.710 1088.000 ;
      LAYER Pwell ;
        RECT 6.290 1080.160 2793.710 1083.680 ;
      LAYER Nwell ;
        RECT 6.290 1075.840 2793.710 1080.160 ;
      LAYER Pwell ;
        RECT 6.290 1072.320 2793.710 1075.840 ;
      LAYER Nwell ;
        RECT 6.290 1068.000 2793.710 1072.320 ;
      LAYER Pwell ;
        RECT 6.290 1064.480 2793.710 1068.000 ;
      LAYER Nwell ;
        RECT 6.290 1060.160 2793.710 1064.480 ;
      LAYER Pwell ;
        RECT 6.290 1056.640 2793.710 1060.160 ;
      LAYER Nwell ;
        RECT 6.290 1052.320 2793.710 1056.640 ;
      LAYER Pwell ;
        RECT 6.290 1048.800 2793.710 1052.320 ;
      LAYER Nwell ;
        RECT 6.290 1044.480 2793.710 1048.800 ;
      LAYER Pwell ;
        RECT 6.290 1040.960 2793.710 1044.480 ;
      LAYER Nwell ;
        RECT 6.290 1036.640 2793.710 1040.960 ;
      LAYER Pwell ;
        RECT 6.290 1033.120 2793.710 1036.640 ;
      LAYER Nwell ;
        RECT 6.290 1028.800 2793.710 1033.120 ;
      LAYER Pwell ;
        RECT 6.290 1025.280 2793.710 1028.800 ;
      LAYER Nwell ;
        RECT 6.290 1020.960 2793.710 1025.280 ;
      LAYER Pwell ;
        RECT 6.290 1017.440 2793.710 1020.960 ;
      LAYER Nwell ;
        RECT 6.290 1013.120 2793.710 1017.440 ;
      LAYER Pwell ;
        RECT 6.290 1009.600 2793.710 1013.120 ;
      LAYER Nwell ;
        RECT 6.290 1005.280 2793.710 1009.600 ;
      LAYER Pwell ;
        RECT 6.290 1001.760 2793.710 1005.280 ;
      LAYER Nwell ;
        RECT 6.290 997.440 2793.710 1001.760 ;
      LAYER Pwell ;
        RECT 6.290 993.920 2793.710 997.440 ;
      LAYER Nwell ;
        RECT 6.290 989.600 2793.710 993.920 ;
      LAYER Pwell ;
        RECT 6.290 986.080 2793.710 989.600 ;
      LAYER Nwell ;
        RECT 6.290 981.760 2793.710 986.080 ;
      LAYER Pwell ;
        RECT 6.290 978.240 2793.710 981.760 ;
      LAYER Nwell ;
        RECT 6.290 973.920 2793.710 978.240 ;
      LAYER Pwell ;
        RECT 6.290 970.400 2793.710 973.920 ;
      LAYER Nwell ;
        RECT 6.290 966.080 2793.710 970.400 ;
      LAYER Pwell ;
        RECT 6.290 962.560 2793.710 966.080 ;
      LAYER Nwell ;
        RECT 6.290 958.240 2793.710 962.560 ;
      LAYER Pwell ;
        RECT 6.290 954.720 2793.710 958.240 ;
      LAYER Nwell ;
        RECT 6.290 950.400 2793.710 954.720 ;
      LAYER Pwell ;
        RECT 6.290 946.880 2793.710 950.400 ;
      LAYER Nwell ;
        RECT 6.290 942.560 2793.710 946.880 ;
      LAYER Pwell ;
        RECT 6.290 939.040 2793.710 942.560 ;
      LAYER Nwell ;
        RECT 6.290 934.720 2793.710 939.040 ;
      LAYER Pwell ;
        RECT 6.290 931.200 2793.710 934.720 ;
      LAYER Nwell ;
        RECT 6.290 926.880 2793.710 931.200 ;
      LAYER Pwell ;
        RECT 6.290 923.360 2793.710 926.880 ;
      LAYER Nwell ;
        RECT 6.290 919.040 2793.710 923.360 ;
      LAYER Pwell ;
        RECT 6.290 915.520 2793.710 919.040 ;
      LAYER Nwell ;
        RECT 6.290 911.200 2793.710 915.520 ;
      LAYER Pwell ;
        RECT 6.290 907.680 2793.710 911.200 ;
      LAYER Nwell ;
        RECT 6.290 903.360 2793.710 907.680 ;
      LAYER Pwell ;
        RECT 6.290 899.840 2793.710 903.360 ;
      LAYER Nwell ;
        RECT 6.290 895.520 2793.710 899.840 ;
      LAYER Pwell ;
        RECT 6.290 892.000 2793.710 895.520 ;
      LAYER Nwell ;
        RECT 6.290 887.680 2793.710 892.000 ;
      LAYER Pwell ;
        RECT 6.290 884.160 2793.710 887.680 ;
      LAYER Nwell ;
        RECT 6.290 879.840 2793.710 884.160 ;
      LAYER Pwell ;
        RECT 6.290 876.320 2793.710 879.840 ;
      LAYER Nwell ;
        RECT 6.290 872.000 2793.710 876.320 ;
      LAYER Pwell ;
        RECT 6.290 868.480 2793.710 872.000 ;
      LAYER Nwell ;
        RECT 6.290 864.160 2793.710 868.480 ;
      LAYER Pwell ;
        RECT 6.290 860.640 2793.710 864.160 ;
      LAYER Nwell ;
        RECT 6.290 856.320 2793.710 860.640 ;
      LAYER Pwell ;
        RECT 6.290 852.800 2793.710 856.320 ;
      LAYER Nwell ;
        RECT 6.290 848.480 2793.710 852.800 ;
      LAYER Pwell ;
        RECT 6.290 844.960 2793.710 848.480 ;
      LAYER Nwell ;
        RECT 6.290 840.640 2793.710 844.960 ;
      LAYER Pwell ;
        RECT 6.290 837.120 2793.710 840.640 ;
      LAYER Nwell ;
        RECT 6.290 832.800 2793.710 837.120 ;
      LAYER Pwell ;
        RECT 6.290 829.280 2793.710 832.800 ;
      LAYER Nwell ;
        RECT 6.290 824.960 2793.710 829.280 ;
      LAYER Pwell ;
        RECT 6.290 821.440 2793.710 824.960 ;
      LAYER Nwell ;
        RECT 6.290 817.120 2793.710 821.440 ;
      LAYER Pwell ;
        RECT 6.290 813.600 2793.710 817.120 ;
      LAYER Nwell ;
        RECT 6.290 809.280 2793.710 813.600 ;
      LAYER Pwell ;
        RECT 6.290 805.760 2793.710 809.280 ;
      LAYER Nwell ;
        RECT 6.290 801.440 2793.710 805.760 ;
      LAYER Pwell ;
        RECT 6.290 797.920 2793.710 801.440 ;
      LAYER Nwell ;
        RECT 6.290 793.600 2793.710 797.920 ;
      LAYER Pwell ;
        RECT 6.290 790.080 2793.710 793.600 ;
      LAYER Nwell ;
        RECT 6.290 785.760 2793.710 790.080 ;
      LAYER Pwell ;
        RECT 6.290 782.240 2793.710 785.760 ;
      LAYER Nwell ;
        RECT 6.290 777.920 2793.710 782.240 ;
      LAYER Pwell ;
        RECT 6.290 774.400 2793.710 777.920 ;
      LAYER Nwell ;
        RECT 6.290 770.080 2793.710 774.400 ;
      LAYER Pwell ;
        RECT 6.290 766.560 2793.710 770.080 ;
      LAYER Nwell ;
        RECT 6.290 762.240 2793.710 766.560 ;
      LAYER Pwell ;
        RECT 6.290 758.720 2793.710 762.240 ;
      LAYER Nwell ;
        RECT 6.290 754.400 2793.710 758.720 ;
      LAYER Pwell ;
        RECT 6.290 750.880 2793.710 754.400 ;
      LAYER Nwell ;
        RECT 6.290 746.560 2793.710 750.880 ;
      LAYER Pwell ;
        RECT 6.290 743.040 2793.710 746.560 ;
      LAYER Nwell ;
        RECT 6.290 738.720 2793.710 743.040 ;
      LAYER Pwell ;
        RECT 6.290 735.200 2793.710 738.720 ;
      LAYER Nwell ;
        RECT 6.290 730.880 2793.710 735.200 ;
      LAYER Pwell ;
        RECT 6.290 727.360 2793.710 730.880 ;
      LAYER Nwell ;
        RECT 6.290 723.040 2793.710 727.360 ;
      LAYER Pwell ;
        RECT 6.290 719.520 2793.710 723.040 ;
      LAYER Nwell ;
        RECT 6.290 715.200 2793.710 719.520 ;
      LAYER Pwell ;
        RECT 6.290 711.680 2793.710 715.200 ;
      LAYER Nwell ;
        RECT 6.290 707.360 2793.710 711.680 ;
      LAYER Pwell ;
        RECT 6.290 703.840 2793.710 707.360 ;
      LAYER Nwell ;
        RECT 6.290 699.520 2793.710 703.840 ;
      LAYER Pwell ;
        RECT 6.290 696.000 2793.710 699.520 ;
      LAYER Nwell ;
        RECT 6.290 691.680 2793.710 696.000 ;
      LAYER Pwell ;
        RECT 6.290 688.160 2793.710 691.680 ;
      LAYER Nwell ;
        RECT 6.290 683.840 2793.710 688.160 ;
      LAYER Pwell ;
        RECT 6.290 680.320 2793.710 683.840 ;
      LAYER Nwell ;
        RECT 6.290 676.000 2793.710 680.320 ;
      LAYER Pwell ;
        RECT 6.290 672.480 2793.710 676.000 ;
      LAYER Nwell ;
        RECT 6.290 668.160 2793.710 672.480 ;
      LAYER Pwell ;
        RECT 6.290 664.640 2793.710 668.160 ;
      LAYER Nwell ;
        RECT 6.290 660.320 2793.710 664.640 ;
      LAYER Pwell ;
        RECT 6.290 656.800 2793.710 660.320 ;
      LAYER Nwell ;
        RECT 6.290 652.480 2793.710 656.800 ;
      LAYER Pwell ;
        RECT 6.290 648.960 2793.710 652.480 ;
      LAYER Nwell ;
        RECT 6.290 644.640 2793.710 648.960 ;
      LAYER Pwell ;
        RECT 6.290 641.120 2793.710 644.640 ;
      LAYER Nwell ;
        RECT 6.290 636.800 2793.710 641.120 ;
      LAYER Pwell ;
        RECT 6.290 633.280 2793.710 636.800 ;
      LAYER Nwell ;
        RECT 6.290 628.960 2793.710 633.280 ;
      LAYER Pwell ;
        RECT 6.290 625.440 2793.710 628.960 ;
      LAYER Nwell ;
        RECT 6.290 621.120 2793.710 625.440 ;
      LAYER Pwell ;
        RECT 6.290 617.600 2793.710 621.120 ;
      LAYER Nwell ;
        RECT 6.290 613.280 2793.710 617.600 ;
      LAYER Pwell ;
        RECT 6.290 609.760 2793.710 613.280 ;
      LAYER Nwell ;
        RECT 6.290 605.440 2793.710 609.760 ;
      LAYER Pwell ;
        RECT 6.290 601.920 2793.710 605.440 ;
      LAYER Nwell ;
        RECT 6.290 597.600 2793.710 601.920 ;
      LAYER Pwell ;
        RECT 6.290 594.080 2793.710 597.600 ;
      LAYER Nwell ;
        RECT 6.290 589.760 2793.710 594.080 ;
      LAYER Pwell ;
        RECT 6.290 586.240 2793.710 589.760 ;
      LAYER Nwell ;
        RECT 6.290 581.920 2793.710 586.240 ;
      LAYER Pwell ;
        RECT 6.290 578.400 2793.710 581.920 ;
      LAYER Nwell ;
        RECT 6.290 574.080 2793.710 578.400 ;
      LAYER Pwell ;
        RECT 6.290 570.560 2793.710 574.080 ;
      LAYER Nwell ;
        RECT 6.290 566.240 2793.710 570.560 ;
      LAYER Pwell ;
        RECT 6.290 562.720 2793.710 566.240 ;
      LAYER Nwell ;
        RECT 6.290 558.400 2793.710 562.720 ;
      LAYER Pwell ;
        RECT 6.290 554.880 2793.710 558.400 ;
      LAYER Nwell ;
        RECT 6.290 550.560 2793.710 554.880 ;
      LAYER Pwell ;
        RECT 6.290 547.040 2793.710 550.560 ;
      LAYER Nwell ;
        RECT 6.290 542.720 2793.710 547.040 ;
      LAYER Pwell ;
        RECT 6.290 539.200 2793.710 542.720 ;
      LAYER Nwell ;
        RECT 6.290 534.880 2793.710 539.200 ;
      LAYER Pwell ;
        RECT 6.290 531.360 2793.710 534.880 ;
      LAYER Nwell ;
        RECT 6.290 527.040 2793.710 531.360 ;
      LAYER Pwell ;
        RECT 6.290 523.520 2793.710 527.040 ;
      LAYER Nwell ;
        RECT 6.290 519.200 2793.710 523.520 ;
      LAYER Pwell ;
        RECT 6.290 515.680 2793.710 519.200 ;
      LAYER Nwell ;
        RECT 6.290 511.360 2793.710 515.680 ;
      LAYER Pwell ;
        RECT 6.290 507.840 2793.710 511.360 ;
      LAYER Nwell ;
        RECT 6.290 503.520 2793.710 507.840 ;
      LAYER Pwell ;
        RECT 6.290 500.000 2793.710 503.520 ;
      LAYER Nwell ;
        RECT 6.290 495.680 2793.710 500.000 ;
      LAYER Pwell ;
        RECT 6.290 492.160 2793.710 495.680 ;
      LAYER Nwell ;
        RECT 6.290 487.840 2793.710 492.160 ;
      LAYER Pwell ;
        RECT 6.290 484.320 2793.710 487.840 ;
      LAYER Nwell ;
        RECT 6.290 480.000 2793.710 484.320 ;
      LAYER Pwell ;
        RECT 6.290 476.480 2793.710 480.000 ;
      LAYER Nwell ;
        RECT 6.290 472.160 2793.710 476.480 ;
      LAYER Pwell ;
        RECT 6.290 468.640 2793.710 472.160 ;
      LAYER Nwell ;
        RECT 6.290 464.320 2793.710 468.640 ;
      LAYER Pwell ;
        RECT 6.290 460.800 2793.710 464.320 ;
      LAYER Nwell ;
        RECT 6.290 456.480 2793.710 460.800 ;
      LAYER Pwell ;
        RECT 6.290 452.960 2793.710 456.480 ;
      LAYER Nwell ;
        RECT 6.290 448.640 2793.710 452.960 ;
      LAYER Pwell ;
        RECT 6.290 445.120 2793.710 448.640 ;
      LAYER Nwell ;
        RECT 6.290 440.800 2793.710 445.120 ;
      LAYER Pwell ;
        RECT 6.290 437.280 2793.710 440.800 ;
      LAYER Nwell ;
        RECT 6.290 432.960 2793.710 437.280 ;
      LAYER Pwell ;
        RECT 6.290 429.440 2793.710 432.960 ;
      LAYER Nwell ;
        RECT 6.290 425.120 2793.710 429.440 ;
      LAYER Pwell ;
        RECT 6.290 421.600 2793.710 425.120 ;
      LAYER Nwell ;
        RECT 6.290 417.280 2793.710 421.600 ;
      LAYER Pwell ;
        RECT 6.290 413.760 2793.710 417.280 ;
      LAYER Nwell ;
        RECT 6.290 409.440 2793.710 413.760 ;
      LAYER Pwell ;
        RECT 6.290 405.920 2793.710 409.440 ;
      LAYER Nwell ;
        RECT 6.290 401.600 2793.710 405.920 ;
      LAYER Pwell ;
        RECT 6.290 398.080 2793.710 401.600 ;
      LAYER Nwell ;
        RECT 6.290 393.760 2793.710 398.080 ;
      LAYER Pwell ;
        RECT 6.290 390.240 2793.710 393.760 ;
      LAYER Nwell ;
        RECT 6.290 385.920 2793.710 390.240 ;
      LAYER Pwell ;
        RECT 6.290 382.400 2793.710 385.920 ;
      LAYER Nwell ;
        RECT 6.290 378.080 2793.710 382.400 ;
      LAYER Pwell ;
        RECT 6.290 374.560 2793.710 378.080 ;
      LAYER Nwell ;
        RECT 6.290 370.240 2793.710 374.560 ;
      LAYER Pwell ;
        RECT 6.290 366.720 2793.710 370.240 ;
      LAYER Nwell ;
        RECT 6.290 362.400 2793.710 366.720 ;
      LAYER Pwell ;
        RECT 6.290 358.880 2793.710 362.400 ;
      LAYER Nwell ;
        RECT 6.290 354.560 2793.710 358.880 ;
      LAYER Pwell ;
        RECT 6.290 351.040 2793.710 354.560 ;
      LAYER Nwell ;
        RECT 6.290 346.720 2793.710 351.040 ;
      LAYER Pwell ;
        RECT 6.290 343.200 2793.710 346.720 ;
      LAYER Nwell ;
        RECT 6.290 338.880 2793.710 343.200 ;
      LAYER Pwell ;
        RECT 6.290 335.360 2793.710 338.880 ;
      LAYER Nwell ;
        RECT 6.290 331.040 2793.710 335.360 ;
      LAYER Pwell ;
        RECT 6.290 327.520 2793.710 331.040 ;
      LAYER Nwell ;
        RECT 6.290 323.200 2793.710 327.520 ;
      LAYER Pwell ;
        RECT 6.290 319.680 2793.710 323.200 ;
      LAYER Nwell ;
        RECT 6.290 315.360 2793.710 319.680 ;
      LAYER Pwell ;
        RECT 6.290 311.840 2793.710 315.360 ;
      LAYER Nwell ;
        RECT 6.290 307.520 2793.710 311.840 ;
      LAYER Pwell ;
        RECT 6.290 304.000 2793.710 307.520 ;
      LAYER Nwell ;
        RECT 6.290 299.680 2793.710 304.000 ;
      LAYER Pwell ;
        RECT 6.290 296.160 2793.710 299.680 ;
      LAYER Nwell ;
        RECT 6.290 291.840 2793.710 296.160 ;
      LAYER Pwell ;
        RECT 6.290 288.320 2793.710 291.840 ;
      LAYER Nwell ;
        RECT 6.290 284.000 2793.710 288.320 ;
      LAYER Pwell ;
        RECT 6.290 280.480 2793.710 284.000 ;
      LAYER Nwell ;
        RECT 6.290 276.160 2793.710 280.480 ;
      LAYER Pwell ;
        RECT 6.290 272.640 2793.710 276.160 ;
      LAYER Nwell ;
        RECT 6.290 268.320 2793.710 272.640 ;
      LAYER Pwell ;
        RECT 6.290 264.800 2793.710 268.320 ;
      LAYER Nwell ;
        RECT 6.290 260.480 2793.710 264.800 ;
      LAYER Pwell ;
        RECT 6.290 256.960 2793.710 260.480 ;
      LAYER Nwell ;
        RECT 6.290 252.640 2793.710 256.960 ;
      LAYER Pwell ;
        RECT 6.290 249.120 2793.710 252.640 ;
      LAYER Nwell ;
        RECT 6.290 244.800 2793.710 249.120 ;
      LAYER Pwell ;
        RECT 6.290 241.280 2793.710 244.800 ;
      LAYER Nwell ;
        RECT 6.290 236.960 2793.710 241.280 ;
      LAYER Pwell ;
        RECT 6.290 233.440 2793.710 236.960 ;
      LAYER Nwell ;
        RECT 6.290 229.120 2793.710 233.440 ;
      LAYER Pwell ;
        RECT 6.290 225.600 2793.710 229.120 ;
      LAYER Nwell ;
        RECT 6.290 221.280 2793.710 225.600 ;
      LAYER Pwell ;
        RECT 6.290 217.760 2793.710 221.280 ;
      LAYER Nwell ;
        RECT 6.290 213.440 2793.710 217.760 ;
      LAYER Pwell ;
        RECT 6.290 209.920 2793.710 213.440 ;
      LAYER Nwell ;
        RECT 6.290 205.600 2793.710 209.920 ;
      LAYER Pwell ;
        RECT 6.290 202.080 2793.710 205.600 ;
      LAYER Nwell ;
        RECT 6.290 197.760 2793.710 202.080 ;
      LAYER Pwell ;
        RECT 6.290 194.240 2793.710 197.760 ;
      LAYER Nwell ;
        RECT 6.290 189.920 2793.710 194.240 ;
      LAYER Pwell ;
        RECT 6.290 186.400 2793.710 189.920 ;
      LAYER Nwell ;
        RECT 6.290 182.080 2793.710 186.400 ;
      LAYER Pwell ;
        RECT 6.290 178.560 2793.710 182.080 ;
      LAYER Nwell ;
        RECT 6.290 174.240 2793.710 178.560 ;
      LAYER Pwell ;
        RECT 6.290 170.720 2793.710 174.240 ;
      LAYER Nwell ;
        RECT 6.290 166.400 2793.710 170.720 ;
      LAYER Pwell ;
        RECT 6.290 162.880 2793.710 166.400 ;
      LAYER Nwell ;
        RECT 6.290 158.560 2793.710 162.880 ;
      LAYER Pwell ;
        RECT 6.290 155.040 2793.710 158.560 ;
      LAYER Nwell ;
        RECT 6.290 150.720 2793.710 155.040 ;
      LAYER Pwell ;
        RECT 6.290 147.200 2793.710 150.720 ;
      LAYER Nwell ;
        RECT 6.290 142.880 2793.710 147.200 ;
      LAYER Pwell ;
        RECT 6.290 139.360 2793.710 142.880 ;
      LAYER Nwell ;
        RECT 6.290 135.040 2793.710 139.360 ;
      LAYER Pwell ;
        RECT 6.290 131.520 2793.710 135.040 ;
      LAYER Nwell ;
        RECT 6.290 127.200 2793.710 131.520 ;
      LAYER Pwell ;
        RECT 6.290 123.680 2793.710 127.200 ;
      LAYER Nwell ;
        RECT 6.290 119.360 2793.710 123.680 ;
      LAYER Pwell ;
        RECT 6.290 115.840 2793.710 119.360 ;
      LAYER Nwell ;
        RECT 6.290 111.520 2793.710 115.840 ;
      LAYER Pwell ;
        RECT 6.290 108.000 2793.710 111.520 ;
      LAYER Nwell ;
        RECT 6.290 103.680 2793.710 108.000 ;
      LAYER Pwell ;
        RECT 6.290 100.160 2793.710 103.680 ;
      LAYER Nwell ;
        RECT 6.290 95.840 2793.710 100.160 ;
      LAYER Pwell ;
        RECT 6.290 92.320 2793.710 95.840 ;
      LAYER Nwell ;
        RECT 6.290 88.000 2793.710 92.320 ;
      LAYER Pwell ;
        RECT 6.290 84.480 2793.710 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 2793.710 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 2793.710 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 2793.710 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 2793.710 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 2793.710 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 2793.710 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 2793.710 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 2793.710 56.640 ;
      LAYER Nwell ;
        RECT 6.290 48.800 2793.710 53.120 ;
      LAYER Pwell ;
        RECT 6.290 45.280 2793.710 48.800 ;
      LAYER Nwell ;
        RECT 6.290 40.960 2793.710 45.280 ;
      LAYER Pwell ;
        RECT 6.290 37.440 2793.710 40.960 ;
      LAYER Nwell ;
        RECT 6.290 33.120 2793.710 37.440 ;
      LAYER Pwell ;
        RECT 6.290 29.600 2793.710 33.120 ;
      LAYER Nwell ;
        RECT 6.290 25.280 2793.710 29.600 ;
      LAYER Pwell ;
        RECT 6.290 21.760 2793.710 25.280 ;
      LAYER Nwell ;
        RECT 6.290 17.440 2793.710 21.760 ;
      LAYER Pwell ;
        RECT 6.290 15.250 2793.710 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 8.550 2793.280 1740.780 ;
      LAYER Metal2 ;
        RECT 22.380 4.300 2788.500 1740.670 ;
        RECT 22.380 4.000 101.620 4.300 ;
        RECT 102.780 4.000 115.060 4.300 ;
        RECT 116.220 4.000 128.500 4.300 ;
        RECT 129.660 4.000 141.940 4.300 ;
        RECT 143.100 4.000 155.380 4.300 ;
        RECT 156.540 4.000 168.820 4.300 ;
        RECT 169.980 4.000 182.260 4.300 ;
        RECT 183.420 4.000 195.700 4.300 ;
        RECT 196.860 4.000 209.140 4.300 ;
        RECT 210.300 4.000 222.580 4.300 ;
        RECT 223.740 4.000 236.020 4.300 ;
        RECT 237.180 4.000 249.460 4.300 ;
        RECT 250.620 4.000 262.900 4.300 ;
        RECT 264.060 4.000 276.340 4.300 ;
        RECT 277.500 4.000 289.780 4.300 ;
        RECT 290.940 4.000 303.220 4.300 ;
        RECT 304.380 4.000 316.660 4.300 ;
        RECT 317.820 4.000 330.100 4.300 ;
        RECT 331.260 4.000 343.540 4.300 ;
        RECT 344.700 4.000 356.980 4.300 ;
        RECT 358.140 4.000 370.420 4.300 ;
        RECT 371.580 4.000 383.860 4.300 ;
        RECT 385.020 4.000 397.300 4.300 ;
        RECT 398.460 4.000 410.740 4.300 ;
        RECT 411.900 4.000 424.180 4.300 ;
        RECT 425.340 4.000 437.620 4.300 ;
        RECT 438.780 4.000 451.060 4.300 ;
        RECT 452.220 4.000 464.500 4.300 ;
        RECT 465.660 4.000 477.940 4.300 ;
        RECT 479.100 4.000 491.380 4.300 ;
        RECT 492.540 4.000 504.820 4.300 ;
        RECT 505.980 4.000 518.260 4.300 ;
        RECT 519.420 4.000 531.700 4.300 ;
        RECT 532.860 4.000 545.140 4.300 ;
        RECT 546.300 4.000 558.580 4.300 ;
        RECT 559.740 4.000 572.020 4.300 ;
        RECT 573.180 4.000 585.460 4.300 ;
        RECT 586.620 4.000 598.900 4.300 ;
        RECT 600.060 4.000 612.340 4.300 ;
        RECT 613.500 4.000 625.780 4.300 ;
        RECT 626.940 4.000 639.220 4.300 ;
        RECT 640.380 4.000 652.660 4.300 ;
        RECT 653.820 4.000 666.100 4.300 ;
        RECT 667.260 4.000 679.540 4.300 ;
        RECT 680.700 4.000 692.980 4.300 ;
        RECT 694.140 4.000 706.420 4.300 ;
        RECT 707.580 4.000 719.860 4.300 ;
        RECT 721.020 4.000 733.300 4.300 ;
        RECT 734.460 4.000 746.740 4.300 ;
        RECT 747.900 4.000 760.180 4.300 ;
        RECT 761.340 4.000 773.620 4.300 ;
        RECT 774.780 4.000 787.060 4.300 ;
        RECT 788.220 4.000 800.500 4.300 ;
        RECT 801.660 4.000 813.940 4.300 ;
        RECT 815.100 4.000 827.380 4.300 ;
        RECT 828.540 4.000 840.820 4.300 ;
        RECT 841.980 4.000 854.260 4.300 ;
        RECT 855.420 4.000 867.700 4.300 ;
        RECT 868.860 4.000 881.140 4.300 ;
        RECT 882.300 4.000 894.580 4.300 ;
        RECT 895.740 4.000 908.020 4.300 ;
        RECT 909.180 4.000 921.460 4.300 ;
        RECT 922.620 4.000 934.900 4.300 ;
        RECT 936.060 4.000 948.340 4.300 ;
        RECT 949.500 4.000 961.780 4.300 ;
        RECT 962.940 4.000 975.220 4.300 ;
        RECT 976.380 4.000 988.660 4.300 ;
        RECT 989.820 4.000 1002.100 4.300 ;
        RECT 1003.260 4.000 1015.540 4.300 ;
        RECT 1016.700 4.000 1028.980 4.300 ;
        RECT 1030.140 4.000 1042.420 4.300 ;
        RECT 1043.580 4.000 1055.860 4.300 ;
        RECT 1057.020 4.000 1069.300 4.300 ;
        RECT 1070.460 4.000 1082.740 4.300 ;
        RECT 1083.900 4.000 1096.180 4.300 ;
        RECT 1097.340 4.000 1109.620 4.300 ;
        RECT 1110.780 4.000 1123.060 4.300 ;
        RECT 1124.220 4.000 1136.500 4.300 ;
        RECT 1137.660 4.000 1149.940 4.300 ;
        RECT 1151.100 4.000 1163.380 4.300 ;
        RECT 1164.540 4.000 1176.820 4.300 ;
        RECT 1177.980 4.000 1190.260 4.300 ;
        RECT 1191.420 4.000 1203.700 4.300 ;
        RECT 1204.860 4.000 1217.140 4.300 ;
        RECT 1218.300 4.000 1230.580 4.300 ;
        RECT 1231.740 4.000 1244.020 4.300 ;
        RECT 1245.180 4.000 1257.460 4.300 ;
        RECT 1258.620 4.000 1270.900 4.300 ;
        RECT 1272.060 4.000 1284.340 4.300 ;
        RECT 1285.500 4.000 1297.780 4.300 ;
        RECT 1298.940 4.000 1311.220 4.300 ;
        RECT 1312.380 4.000 1324.660 4.300 ;
        RECT 1325.820 4.000 1338.100 4.300 ;
        RECT 1339.260 4.000 1351.540 4.300 ;
        RECT 1352.700 4.000 1364.980 4.300 ;
        RECT 1366.140 4.000 1378.420 4.300 ;
        RECT 1379.580 4.000 1391.860 4.300 ;
        RECT 1393.020 4.000 1405.300 4.300 ;
        RECT 1406.460 4.000 1418.740 4.300 ;
        RECT 1419.900 4.000 1432.180 4.300 ;
        RECT 1433.340 4.000 1445.620 4.300 ;
        RECT 1446.780 4.000 1459.060 4.300 ;
        RECT 1460.220 4.000 1472.500 4.300 ;
        RECT 1473.660 4.000 1485.940 4.300 ;
        RECT 1487.100 4.000 1499.380 4.300 ;
        RECT 1500.540 4.000 1512.820 4.300 ;
        RECT 1513.980 4.000 1526.260 4.300 ;
        RECT 1527.420 4.000 1539.700 4.300 ;
        RECT 1540.860 4.000 1553.140 4.300 ;
        RECT 1554.300 4.000 1566.580 4.300 ;
        RECT 1567.740 4.000 1580.020 4.300 ;
        RECT 1581.180 4.000 1593.460 4.300 ;
        RECT 1594.620 4.000 1606.900 4.300 ;
        RECT 1608.060 4.000 1620.340 4.300 ;
        RECT 1621.500 4.000 1633.780 4.300 ;
        RECT 1634.940 4.000 1647.220 4.300 ;
        RECT 1648.380 4.000 1660.660 4.300 ;
        RECT 1661.820 4.000 1674.100 4.300 ;
        RECT 1675.260 4.000 1687.540 4.300 ;
        RECT 1688.700 4.000 1700.980 4.300 ;
        RECT 1702.140 4.000 1714.420 4.300 ;
        RECT 1715.580 4.000 1727.860 4.300 ;
        RECT 1729.020 4.000 1741.300 4.300 ;
        RECT 1742.460 4.000 1754.740 4.300 ;
        RECT 1755.900 4.000 1768.180 4.300 ;
        RECT 1769.340 4.000 1781.620 4.300 ;
        RECT 1782.780 4.000 1795.060 4.300 ;
        RECT 1796.220 4.000 1808.500 4.300 ;
        RECT 1809.660 4.000 1821.940 4.300 ;
        RECT 1823.100 4.000 1835.380 4.300 ;
        RECT 1836.540 4.000 1848.820 4.300 ;
        RECT 1849.980 4.000 1862.260 4.300 ;
        RECT 1863.420 4.000 1875.700 4.300 ;
        RECT 1876.860 4.000 1889.140 4.300 ;
        RECT 1890.300 4.000 1902.580 4.300 ;
        RECT 1903.740 4.000 1916.020 4.300 ;
        RECT 1917.180 4.000 1929.460 4.300 ;
        RECT 1930.620 4.000 1942.900 4.300 ;
        RECT 1944.060 4.000 1956.340 4.300 ;
        RECT 1957.500 4.000 1969.780 4.300 ;
        RECT 1970.940 4.000 1983.220 4.300 ;
        RECT 1984.380 4.000 1996.660 4.300 ;
        RECT 1997.820 4.000 2010.100 4.300 ;
        RECT 2011.260 4.000 2023.540 4.300 ;
        RECT 2024.700 4.000 2036.980 4.300 ;
        RECT 2038.140 4.000 2050.420 4.300 ;
        RECT 2051.580 4.000 2063.860 4.300 ;
        RECT 2065.020 4.000 2077.300 4.300 ;
        RECT 2078.460 4.000 2090.740 4.300 ;
        RECT 2091.900 4.000 2104.180 4.300 ;
        RECT 2105.340 4.000 2117.620 4.300 ;
        RECT 2118.780 4.000 2131.060 4.300 ;
        RECT 2132.220 4.000 2144.500 4.300 ;
        RECT 2145.660 4.000 2157.940 4.300 ;
        RECT 2159.100 4.000 2171.380 4.300 ;
        RECT 2172.540 4.000 2184.820 4.300 ;
        RECT 2185.980 4.000 2198.260 4.300 ;
        RECT 2199.420 4.000 2211.700 4.300 ;
        RECT 2212.860 4.000 2225.140 4.300 ;
        RECT 2226.300 4.000 2238.580 4.300 ;
        RECT 2239.740 4.000 2252.020 4.300 ;
        RECT 2253.180 4.000 2265.460 4.300 ;
        RECT 2266.620 4.000 2278.900 4.300 ;
        RECT 2280.060 4.000 2292.340 4.300 ;
        RECT 2293.500 4.000 2305.780 4.300 ;
        RECT 2306.940 4.000 2319.220 4.300 ;
        RECT 2320.380 4.000 2332.660 4.300 ;
        RECT 2333.820 4.000 2346.100 4.300 ;
        RECT 2347.260 4.000 2359.540 4.300 ;
        RECT 2360.700 4.000 2372.980 4.300 ;
        RECT 2374.140 4.000 2386.420 4.300 ;
        RECT 2387.580 4.000 2399.860 4.300 ;
        RECT 2401.020 4.000 2413.300 4.300 ;
        RECT 2414.460 4.000 2426.740 4.300 ;
        RECT 2427.900 4.000 2440.180 4.300 ;
        RECT 2441.340 4.000 2453.620 4.300 ;
        RECT 2454.780 4.000 2467.060 4.300 ;
        RECT 2468.220 4.000 2480.500 4.300 ;
        RECT 2481.660 4.000 2493.940 4.300 ;
        RECT 2495.100 4.000 2507.380 4.300 ;
        RECT 2508.540 4.000 2520.820 4.300 ;
        RECT 2521.980 4.000 2534.260 4.300 ;
        RECT 2535.420 4.000 2547.700 4.300 ;
        RECT 2548.860 4.000 2561.140 4.300 ;
        RECT 2562.300 4.000 2574.580 4.300 ;
        RECT 2575.740 4.000 2588.020 4.300 ;
        RECT 2589.180 4.000 2601.460 4.300 ;
        RECT 2602.620 4.000 2614.900 4.300 ;
        RECT 2616.060 4.000 2628.340 4.300 ;
        RECT 2629.500 4.000 2641.780 4.300 ;
        RECT 2642.940 4.000 2655.220 4.300 ;
        RECT 2656.380 4.000 2668.660 4.300 ;
        RECT 2669.820 4.000 2682.100 4.300 ;
        RECT 2683.260 4.000 2695.540 4.300 ;
        RECT 2696.700 4.000 2788.500 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 15.540 2788.550 1740.620 ;
  END
END user_proj_example
END LIBRARY

